`define FONT_HEIGHT 16
`define FONT_WIDTH  8

module font_vt323_8x16
#(
  parameter XY_BIT_DEPTH = 8
)
(
  input wire  [XY_BIT_DEPTH-1:0] sym_x,
  input wire  [XY_BIT_DEPTH-1:0] sym_y,
  input wire  [7:0]              sym_code,
  output wire                    sym_pixel
);

  wire [`FONT_WIDTH-1:0] font [`FONT_HEIGHT-1:0] [255:0];

// Here all font bits should be assigned
	assign font[0][0] = 8'b11111111;
	assign font[1][0] = 8'b11111111;
	assign font[2][0] = 8'b11111111;
	assign font[3][0] = 8'b11111111;
	assign font[4][0] = 8'b11111111;
	assign font[5][0] = 8'b11111111;
	assign font[6][0] = 8'b11111111;
	assign font[7][0] = 8'b11111111;
	assign font[8][0] = 8'b11111111;
	assign font[9][0] = 8'b11111111;
	assign font[10][0] = 8'b11111111;
	assign font[11][0] = 8'b11111111;
	assign font[12][0] = 8'b11111111;
	assign font[13][0] = 8'b11111111;
	assign font[14][0] = 8'b11111111;
	assign font[15][0] = 8'b11111111;

	assign font[0][1] = 8'b11111111;
	assign font[1][1] = 8'b11111111;
	assign font[2][1] = 8'b11111111;
	assign font[3][1] = 8'b11111111;
	assign font[4][1] = 8'b11111111;
	assign font[5][1] = 8'b11111111;
	assign font[6][1] = 8'b11111111;
	assign font[7][1] = 8'b11111111;
	assign font[8][1] = 8'b11111111;
	assign font[9][1] = 8'b11111111;
	assign font[10][1] = 8'b11111111;
	assign font[11][1] = 8'b11111111;
	assign font[12][1] = 8'b11111111;
	assign font[13][1] = 8'b11111111;
	assign font[14][1] = 8'b11111111;
	assign font[15][1] = 8'b11111111;

	assign font[0][2] = 8'b11111111;
	assign font[1][2] = 8'b11111111;
	assign font[2][2] = 8'b11111111;
	assign font[3][2] = 8'b11111111;
	assign font[4][2] = 8'b11111111;
	assign font[5][2] = 8'b11111111;
	assign font[6][2] = 8'b11111111;
	assign font[7][2] = 8'b11111111;
	assign font[8][2] = 8'b11111111;
	assign font[9][2] = 8'b11111111;
	assign font[10][2] = 8'b11111111;
	assign font[11][2] = 8'b11111111;
	assign font[12][2] = 8'b11111111;
	assign font[13][2] = 8'b11111111;
	assign font[14][2] = 8'b11111111;
	assign font[15][2] = 8'b11111111;

	assign font[0][3] = 8'b11111111;
	assign font[1][3] = 8'b11111111;
	assign font[2][3] = 8'b11111111;
	assign font[3][3] = 8'b11111111;
	assign font[4][3] = 8'b11111111;
	assign font[5][3] = 8'b11111111;
	assign font[6][3] = 8'b11111111;
	assign font[7][3] = 8'b11111111;
	assign font[8][3] = 8'b11111111;
	assign font[9][3] = 8'b11111111;
	assign font[10][3] = 8'b11111111;
	assign font[11][3] = 8'b11111111;
	assign font[12][3] = 8'b11111111;
	assign font[13][3] = 8'b11111111;
	assign font[14][3] = 8'b11111111;
	assign font[15][3] = 8'b11111111;

	assign font[0][4] = 8'b11111111;
	assign font[1][4] = 8'b11111111;
	assign font[2][4] = 8'b11111111;
	assign font[3][4] = 8'b11111111;
	assign font[4][4] = 8'b11111111;
	assign font[5][4] = 8'b11111111;
	assign font[6][4] = 8'b11111111;
	assign font[7][4] = 8'b11111111;
	assign font[8][4] = 8'b11111111;
	assign font[9][4] = 8'b11111111;
	assign font[10][4] = 8'b11111111;
	assign font[11][4] = 8'b11111111;
	assign font[12][4] = 8'b11111111;
	assign font[13][4] = 8'b11111111;
	assign font[14][4] = 8'b11111111;
	assign font[15][4] = 8'b11111111;

	assign font[0][5] = 8'b11111111;
	assign font[1][5] = 8'b11111111;
	assign font[2][5] = 8'b11111111;
	assign font[3][5] = 8'b11111111;
	assign font[4][5] = 8'b11111111;
	assign font[5][5] = 8'b11111111;
	assign font[6][5] = 8'b11111111;
	assign font[7][5] = 8'b11111111;
	assign font[8][5] = 8'b11111111;
	assign font[9][5] = 8'b11111111;
	assign font[10][5] = 8'b11111111;
	assign font[11][5] = 8'b11111111;
	assign font[12][5] = 8'b11111111;
	assign font[13][5] = 8'b11111111;
	assign font[14][5] = 8'b11111111;
	assign font[15][5] = 8'b11111111;

	assign font[0][6] = 8'b11111111;
	assign font[1][6] = 8'b11111111;
	assign font[2][6] = 8'b11111111;
	assign font[3][6] = 8'b11111111;
	assign font[4][6] = 8'b11111111;
	assign font[5][6] = 8'b11111111;
	assign font[6][6] = 8'b11111111;
	assign font[7][6] = 8'b11111111;
	assign font[8][6] = 8'b11111111;
	assign font[9][6] = 8'b11111111;
	assign font[10][6] = 8'b11111111;
	assign font[11][6] = 8'b11111111;
	assign font[12][6] = 8'b11111111;
	assign font[13][6] = 8'b11111111;
	assign font[14][6] = 8'b11111111;
	assign font[15][6] = 8'b11111111;

	assign font[0][7] = 8'b11111111;
	assign font[1][7] = 8'b11111111;
	assign font[2][7] = 8'b11111111;
	assign font[3][7] = 8'b11111111;
	assign font[4][7] = 8'b11111111;
	assign font[5][7] = 8'b11111111;
	assign font[6][7] = 8'b11111111;
	assign font[7][7] = 8'b11111111;
	assign font[8][7] = 8'b11111111;
	assign font[9][7] = 8'b11111111;
	assign font[10][7] = 8'b11111111;
	assign font[11][7] = 8'b11111111;
	assign font[12][7] = 8'b11111111;
	assign font[13][7] = 8'b11111111;
	assign font[14][7] = 8'b11111111;
	assign font[15][7] = 8'b11111111;

	assign font[0][8] = 8'b11111111;
	assign font[1][8] = 8'b11111111;
	assign font[2][8] = 8'b11111111;
	assign font[3][8] = 8'b11111111;
	assign font[4][8] = 8'b11111111;
	assign font[5][8] = 8'b11111111;
	assign font[6][8] = 8'b11111111;
	assign font[7][8] = 8'b11111111;
	assign font[8][8] = 8'b11111111;
	assign font[9][8] = 8'b11111111;
	assign font[10][8] = 8'b11111111;
	assign font[11][8] = 8'b11111111;
	assign font[12][8] = 8'b11111111;
	assign font[13][8] = 8'b11111111;
	assign font[14][8] = 8'b11111111;
	assign font[15][8] = 8'b11111111;

	assign font[0][9] = 8'b11111111;
	assign font[1][9] = 8'b11111111;
	assign font[2][9] = 8'b11111111;
	assign font[3][9] = 8'b11111111;
	assign font[4][9] = 8'b11111111;
	assign font[5][9] = 8'b11111111;
	assign font[6][9] = 8'b11111111;
	assign font[7][9] = 8'b11111111;
	assign font[8][9] = 8'b11111111;
	assign font[9][9] = 8'b11111111;
	assign font[10][9] = 8'b11111111;
	assign font[11][9] = 8'b11111111;
	assign font[12][9] = 8'b11111111;
	assign font[13][9] = 8'b11111111;
	assign font[14][9] = 8'b11111111;
	assign font[15][9] = 8'b11111111;

	assign font[0][10] = 8'b11111111;
	assign font[1][10] = 8'b11111111;
	assign font[2][10] = 8'b11111111;
	assign font[3][10] = 8'b11111111;
	assign font[4][10] = 8'b11111111;
	assign font[5][10] = 8'b11111111;
	assign font[6][10] = 8'b11111111;
	assign font[7][10] = 8'b11111111;
	assign font[8][10] = 8'b11111111;
	assign font[9][10] = 8'b11111111;
	assign font[10][10] = 8'b11111111;
	assign font[11][10] = 8'b11111111;
	assign font[12][10] = 8'b11111111;
	assign font[13][10] = 8'b11111111;
	assign font[14][10] = 8'b11111111;
	assign font[15][10] = 8'b11111111;

	assign font[0][11] = 8'b11111111;
	assign font[1][11] = 8'b11111111;
	assign font[2][11] = 8'b11111111;
	assign font[3][11] = 8'b11111111;
	assign font[4][11] = 8'b11111111;
	assign font[5][11] = 8'b11111111;
	assign font[6][11] = 8'b11111111;
	assign font[7][11] = 8'b11111111;
	assign font[8][11] = 8'b11111111;
	assign font[9][11] = 8'b11111111;
	assign font[10][11] = 8'b11111111;
	assign font[11][11] = 8'b11111111;
	assign font[12][11] = 8'b11111111;
	assign font[13][11] = 8'b11111111;
	assign font[14][11] = 8'b11111111;
	assign font[15][11] = 8'b11111111;

	assign font[0][12] = 8'b11111111;
	assign font[1][12] = 8'b11111111;
	assign font[2][12] = 8'b11111111;
	assign font[3][12] = 8'b11111111;
	assign font[4][12] = 8'b11111111;
	assign font[5][12] = 8'b11111111;
	assign font[6][12] = 8'b11111111;
	assign font[7][12] = 8'b11111111;
	assign font[8][12] = 8'b11111111;
	assign font[9][12] = 8'b11111111;
	assign font[10][12] = 8'b11111111;
	assign font[11][12] = 8'b11111111;
	assign font[12][12] = 8'b11111111;
	assign font[13][12] = 8'b11111111;
	assign font[14][12] = 8'b11111111;
	assign font[15][12] = 8'b11111111;

	assign font[0][13] = 8'b11111111;
	assign font[1][13] = 8'b11111111;
	assign font[2][13] = 8'b11111111;
	assign font[3][13] = 8'b11111111;
	assign font[4][13] = 8'b11111111;
	assign font[5][13] = 8'b11111111;
	assign font[6][13] = 8'b11111111;
	assign font[7][13] = 8'b11111111;
	assign font[8][13] = 8'b11111111;
	assign font[9][13] = 8'b11111111;
	assign font[10][13] = 8'b11111111;
	assign font[11][13] = 8'b11111111;
	assign font[12][13] = 8'b11111111;
	assign font[13][13] = 8'b11111111;
	assign font[14][13] = 8'b11111111;
	assign font[15][13] = 8'b11111111;

	assign font[0][14] = 8'b11111111;
	assign font[1][14] = 8'b11111111;
	assign font[2][14] = 8'b11111111;
	assign font[3][14] = 8'b11111111;
	assign font[4][14] = 8'b11111111;
	assign font[5][14] = 8'b11111111;
	assign font[6][14] = 8'b11111111;
	assign font[7][14] = 8'b11111111;
	assign font[8][14] = 8'b11111111;
	assign font[9][14] = 8'b11111111;
	assign font[10][14] = 8'b11111111;
	assign font[11][14] = 8'b11111111;
	assign font[12][14] = 8'b11111111;
	assign font[13][14] = 8'b11111111;
	assign font[14][14] = 8'b11111111;
	assign font[15][14] = 8'b11111111;

	assign font[0][15] = 8'b11111111;
	assign font[1][15] = 8'b11111111;
	assign font[2][15] = 8'b11111111;
	assign font[3][15] = 8'b11111111;
	assign font[4][15] = 8'b11111111;
	assign font[5][15] = 8'b11111111;
	assign font[6][15] = 8'b11111111;
	assign font[7][15] = 8'b11111111;
	assign font[8][15] = 8'b11111111;
	assign font[9][15] = 8'b11111111;
	assign font[10][15] = 8'b11111111;
	assign font[11][15] = 8'b11111111;
	assign font[12][15] = 8'b11111111;
	assign font[13][15] = 8'b11111111;
	assign font[14][15] = 8'b11111111;
	assign font[15][15] = 8'b11111111;

	assign font[0][16] = 8'b11111111;
	assign font[1][16] = 8'b11111111;
	assign font[2][16] = 8'b11111111;
	assign font[3][16] = 8'b11111111;
	assign font[4][16] = 8'b11111111;
	assign font[5][16] = 8'b11111111;
	assign font[6][16] = 8'b11111111;
	assign font[7][16] = 8'b11111111;
	assign font[8][16] = 8'b11111111;
	assign font[9][16] = 8'b11111111;
	assign font[10][16] = 8'b11111111;
	assign font[11][16] = 8'b11111111;
	assign font[12][16] = 8'b11111111;
	assign font[13][16] = 8'b11111111;
	assign font[14][16] = 8'b11111111;
	assign font[15][16] = 8'b11111111;

	assign font[0][17] = 8'b11111111;
	assign font[1][17] = 8'b11111111;
	assign font[2][17] = 8'b11111111;
	assign font[3][17] = 8'b11111111;
	assign font[4][17] = 8'b11111111;
	assign font[5][17] = 8'b11111111;
	assign font[6][17] = 8'b11111111;
	assign font[7][17] = 8'b11111111;
	assign font[8][17] = 8'b11111111;
	assign font[9][17] = 8'b11111111;
	assign font[10][17] = 8'b11111111;
	assign font[11][17] = 8'b11111111;
	assign font[12][17] = 8'b11111111;
	assign font[13][17] = 8'b11111111;
	assign font[14][17] = 8'b11111111;
	assign font[15][17] = 8'b11111111;

	assign font[0][18] = 8'b11111111;
	assign font[1][18] = 8'b11111111;
	assign font[2][18] = 8'b11111111;
	assign font[3][18] = 8'b11111111;
	assign font[4][18] = 8'b11111111;
	assign font[5][18] = 8'b11111111;
	assign font[6][18] = 8'b11111111;
	assign font[7][18] = 8'b11111111;
	assign font[8][18] = 8'b11111111;
	assign font[9][18] = 8'b11111111;
	assign font[10][18] = 8'b11111111;
	assign font[11][18] = 8'b11111111;
	assign font[12][18] = 8'b11111111;
	assign font[13][18] = 8'b11111111;
	assign font[14][18] = 8'b11111111;
	assign font[15][18] = 8'b11111111;

	assign font[0][19] = 8'b11111111;
	assign font[1][19] = 8'b11111111;
	assign font[2][19] = 8'b11111111;
	assign font[3][19] = 8'b11111111;
	assign font[4][19] = 8'b11111111;
	assign font[5][19] = 8'b11111111;
	assign font[6][19] = 8'b11111111;
	assign font[7][19] = 8'b11111111;
	assign font[8][19] = 8'b11111111;
	assign font[9][19] = 8'b11111111;
	assign font[10][19] = 8'b11111111;
	assign font[11][19] = 8'b11111111;
	assign font[12][19] = 8'b11111111;
	assign font[13][19] = 8'b11111111;
	assign font[14][19] = 8'b11111111;
	assign font[15][19] = 8'b11111111;

	assign font[0][20] = 8'b11111111;
	assign font[1][20] = 8'b11111111;
	assign font[2][20] = 8'b11111111;
	assign font[3][20] = 8'b11111111;
	assign font[4][20] = 8'b11111111;
	assign font[5][20] = 8'b11111111;
	assign font[6][20] = 8'b11111111;
	assign font[7][20] = 8'b11111111;
	assign font[8][20] = 8'b11111111;
	assign font[9][20] = 8'b11111111;
	assign font[10][20] = 8'b11111111;
	assign font[11][20] = 8'b11111111;
	assign font[12][20] = 8'b11111111;
	assign font[13][20] = 8'b11111111;
	assign font[14][20] = 8'b11111111;
	assign font[15][20] = 8'b11111111;

	assign font[0][21] = 8'b11111111;
	assign font[1][21] = 8'b11111111;
	assign font[2][21] = 8'b11111111;
	assign font[3][21] = 8'b11111111;
	assign font[4][21] = 8'b11111111;
	assign font[5][21] = 8'b11111111;
	assign font[6][21] = 8'b11111111;
	assign font[7][21] = 8'b11111111;
	assign font[8][21] = 8'b11111111;
	assign font[9][21] = 8'b11111111;
	assign font[10][21] = 8'b11111111;
	assign font[11][21] = 8'b11111111;
	assign font[12][21] = 8'b11111111;
	assign font[13][21] = 8'b11111111;
	assign font[14][21] = 8'b11111111;
	assign font[15][21] = 8'b11111111;

	assign font[0][22] = 8'b11111111;
	assign font[1][22] = 8'b11111111;
	assign font[2][22] = 8'b11111111;
	assign font[3][22] = 8'b11111111;
	assign font[4][22] = 8'b11111111;
	assign font[5][22] = 8'b11111111;
	assign font[6][22] = 8'b11111111;
	assign font[7][22] = 8'b11111111;
	assign font[8][22] = 8'b11111111;
	assign font[9][22] = 8'b11111111;
	assign font[10][22] = 8'b11111111;
	assign font[11][22] = 8'b11111111;
	assign font[12][22] = 8'b11111111;
	assign font[13][22] = 8'b11111111;
	assign font[14][22] = 8'b11111111;
	assign font[15][22] = 8'b11111111;

	assign font[0][23] = 8'b11111111;
	assign font[1][23] = 8'b11111111;
	assign font[2][23] = 8'b11111111;
	assign font[3][23] = 8'b11111111;
	assign font[4][23] = 8'b11111111;
	assign font[5][23] = 8'b11111111;
	assign font[6][23] = 8'b11111111;
	assign font[7][23] = 8'b11111111;
	assign font[8][23] = 8'b11111111;
	assign font[9][23] = 8'b11111111;
	assign font[10][23] = 8'b11111111;
	assign font[11][23] = 8'b11111111;
	assign font[12][23] = 8'b11111111;
	assign font[13][23] = 8'b11111111;
	assign font[14][23] = 8'b11111111;
	assign font[15][23] = 8'b11111111;

	assign font[0][24] = 8'b11111111;
	assign font[1][24] = 8'b11111111;
	assign font[2][24] = 8'b11111111;
	assign font[3][24] = 8'b11111111;
	assign font[4][24] = 8'b11111111;
	assign font[5][24] = 8'b11111111;
	assign font[6][24] = 8'b11111111;
	assign font[7][24] = 8'b11111111;
	assign font[8][24] = 8'b11111111;
	assign font[9][24] = 8'b11111111;
	assign font[10][24] = 8'b11111111;
	assign font[11][24] = 8'b11111111;
	assign font[12][24] = 8'b11111111;
	assign font[13][24] = 8'b11111111;
	assign font[14][24] = 8'b11111111;
	assign font[15][24] = 8'b11111111;

	assign font[0][25] = 8'b11111111;
	assign font[1][25] = 8'b11111111;
	assign font[2][25] = 8'b11111111;
	assign font[3][25] = 8'b11111111;
	assign font[4][25] = 8'b11111111;
	assign font[5][25] = 8'b11111111;
	assign font[6][25] = 8'b11111111;
	assign font[7][25] = 8'b11111111;
	assign font[8][25] = 8'b11111111;
	assign font[9][25] = 8'b11111111;
	assign font[10][25] = 8'b11111111;
	assign font[11][25] = 8'b11111111;
	assign font[12][25] = 8'b11111111;
	assign font[13][25] = 8'b11111111;
	assign font[14][25] = 8'b11111111;
	assign font[15][25] = 8'b11111111;

	assign font[0][26] = 8'b11111111;
	assign font[1][26] = 8'b11111111;
	assign font[2][26] = 8'b11111111;
	assign font[3][26] = 8'b11111111;
	assign font[4][26] = 8'b11111111;
	assign font[5][26] = 8'b11111111;
	assign font[6][26] = 8'b11111111;
	assign font[7][26] = 8'b11111111;
	assign font[8][26] = 8'b11111111;
	assign font[9][26] = 8'b11111111;
	assign font[10][26] = 8'b11111111;
	assign font[11][26] = 8'b11111111;
	assign font[12][26] = 8'b11111111;
	assign font[13][26] = 8'b11111111;
	assign font[14][26] = 8'b11111111;
	assign font[15][26] = 8'b11111111;

	assign font[0][27] = 8'b11111111;
	assign font[1][27] = 8'b11111111;
	assign font[2][27] = 8'b11111111;
	assign font[3][27] = 8'b11111111;
	assign font[4][27] = 8'b11111111;
	assign font[5][27] = 8'b11111111;
	assign font[6][27] = 8'b11111111;
	assign font[7][27] = 8'b11111111;
	assign font[8][27] = 8'b11111111;
	assign font[9][27] = 8'b11111111;
	assign font[10][27] = 8'b11111111;
	assign font[11][27] = 8'b11111111;
	assign font[12][27] = 8'b11111111;
	assign font[13][27] = 8'b11111111;
	assign font[14][27] = 8'b11111111;
	assign font[15][27] = 8'b11111111;

	assign font[0][28] = 8'b11111111;
	assign font[1][28] = 8'b11111111;
	assign font[2][28] = 8'b11111111;
	assign font[3][28] = 8'b11111111;
	assign font[4][28] = 8'b11111111;
	assign font[5][28] = 8'b11111111;
	assign font[6][28] = 8'b11111111;
	assign font[7][28] = 8'b11111111;
	assign font[8][28] = 8'b11111111;
	assign font[9][28] = 8'b11111111;
	assign font[10][28] = 8'b11111111;
	assign font[11][28] = 8'b11111111;
	assign font[12][28] = 8'b11111111;
	assign font[13][28] = 8'b11111111;
	assign font[14][28] = 8'b11111111;
	assign font[15][28] = 8'b11111111;

	assign font[0][29] = 8'b11111111;
	assign font[1][29] = 8'b11111111;
	assign font[2][29] = 8'b11111111;
	assign font[3][29] = 8'b11111111;
	assign font[4][29] = 8'b11111111;
	assign font[5][29] = 8'b11111111;
	assign font[6][29] = 8'b11111111;
	assign font[7][29] = 8'b11111111;
	assign font[8][29] = 8'b11111111;
	assign font[9][29] = 8'b11111111;
	assign font[10][29] = 8'b11111111;
	assign font[11][29] = 8'b11111111;
	assign font[12][29] = 8'b11111111;
	assign font[13][29] = 8'b11111111;
	assign font[14][29] = 8'b11111111;
	assign font[15][29] = 8'b11111111;

	assign font[0][30] = 8'b11111111;
	assign font[1][30] = 8'b11111111;
	assign font[2][30] = 8'b11111111;
	assign font[3][30] = 8'b11111111;
	assign font[4][30] = 8'b11111111;
	assign font[5][30] = 8'b11111111;
	assign font[6][30] = 8'b11111111;
	assign font[7][30] = 8'b11111111;
	assign font[8][30] = 8'b11111111;
	assign font[9][30] = 8'b11111111;
	assign font[10][30] = 8'b11111111;
	assign font[11][30] = 8'b11111111;
	assign font[12][30] = 8'b11111111;
	assign font[13][30] = 8'b11111111;
	assign font[14][30] = 8'b11111111;
	assign font[15][30] = 8'b11111111;

	assign font[0][31] = 8'b11111111;
	assign font[1][31] = 8'b11111111;
	assign font[2][31] = 8'b11111111;
	assign font[3][31] = 8'b11111111;
	assign font[4][31] = 8'b11111111;
	assign font[5][31] = 8'b11111111;
	assign font[6][31] = 8'b11111111;
	assign font[7][31] = 8'b11111111;
	assign font[8][31] = 8'b11111111;
	assign font[9][31] = 8'b11111111;
	assign font[10][31] = 8'b11111111;
	assign font[11][31] = 8'b11111111;
	assign font[12][31] = 8'b11111111;
	assign font[13][31] = 8'b11111111;
	assign font[14][31] = 8'b11111111;
	assign font[15][31] = 8'b11111111;

	assign font[0][32] = 8'b11111111;
	assign font[1][32] = 8'b11111111;
	assign font[2][32] = 8'b11111111;
	assign font[3][32] = 8'b11111111;
	assign font[4][32] = 8'b11111111;
	assign font[5][32] = 8'b11111111;
	assign font[6][32] = 8'b11111111;
	assign font[7][32] = 8'b11111111;
	assign font[8][32] = 8'b11111111;
	assign font[9][32] = 8'b11111111;
	assign font[10][32] = 8'b11111111;
	assign font[11][32] = 8'b11111111;
	assign font[12][32] = 8'b11111111;
	assign font[13][32] = 8'b11111111;
	assign font[14][32] = 8'b11111111;
	assign font[15][32] = 8'b11111111;

	assign font[0][33] = 8'b00000000;
	assign font[1][33] = 8'b00000000;
	assign font[2][33] = 8'b00000000;
	assign font[3][33] = 8'b00000000;
	assign font[4][33] = 8'b00010000;
	assign font[5][33] = 8'b00010000;
	assign font[6][33] = 8'b00010000;
	assign font[7][33] = 8'b00010000;
	assign font[8][33] = 8'b00010000;
	assign font[9][33] = 8'b00010000;
	assign font[10][33] = 8'b00000000;
	assign font[11][33] = 8'b00000000;
	assign font[12][33] = 8'b00000000;
	assign font[13][33] = 8'b00010000;
	assign font[14][33] = 8'b00000000;
	assign font[15][33] = 8'b00000000;

	assign font[0][34] = 8'b00000000;
	assign font[1][34] = 8'b00000000;
	assign font[2][34] = 8'b00000000;
	assign font[3][34] = 8'b00000000;
	assign font[4][34] = 8'b00100100;
	assign font[5][34] = 8'b00100100;
	assign font[6][34] = 8'b00000000;
	assign font[7][34] = 8'b00000000;
	assign font[8][34] = 8'b00000000;
	assign font[9][34] = 8'b00000000;
	assign font[10][34] = 8'b00000000;
	assign font[11][34] = 8'b00000000;
	assign font[12][34] = 8'b00000000;
	assign font[13][34] = 8'b00000000;
	assign font[14][34] = 8'b00000000;
	assign font[15][34] = 8'b00000000;

	assign font[0][35] = 8'b00000000;
	assign font[1][35] = 8'b00000000;
	assign font[2][35] = 8'b00000000;
	assign font[3][35] = 8'b00000000;
	assign font[4][35] = 8'b00000000;
	assign font[5][35] = 8'b00000000;
	assign font[6][35] = 8'b00101000;
	assign font[7][35] = 8'b01111100;
	assign font[8][35] = 8'b00101100;
	assign font[9][35] = 8'b00101000;
	assign font[10][35] = 8'b00101000;
	assign font[11][35] = 8'b00101000;
	assign font[12][35] = 8'b01111100;
	assign font[13][35] = 8'b00101000;
	assign font[14][35] = 8'b00000000;
	assign font[15][35] = 8'b00000000;

	assign font[0][36] = 8'b00000000;
	assign font[1][36] = 8'b00000000;
	assign font[2][36] = 8'b00000000;
	assign font[3][36] = 8'b00000000;
	assign font[4][36] = 8'b00010000;
	assign font[5][36] = 8'b00010000;
	assign font[6][36] = 8'b00111000;
	assign font[7][36] = 8'b01010000;
	assign font[8][36] = 8'b01010000;
	assign font[9][36] = 8'b00111000;
	assign font[10][36] = 8'b00010100;
	assign font[11][36] = 8'b00011000;
	assign font[12][36] = 8'b00111000;
	assign font[13][36] = 8'b00010000;
	assign font[14][36] = 8'b00000000;
	assign font[15][36] = 8'b00000000;

	assign font[0][37] = 8'b00000000;
	assign font[1][37] = 8'b00000000;
	assign font[2][37] = 8'b00000000;
	assign font[3][37] = 8'b00000000;
	assign font[4][37] = 8'b01101000;
	assign font[5][37] = 8'b01101000;
	assign font[6][37] = 8'b01101000;
	assign font[7][37] = 8'b01101000;
	assign font[8][37] = 8'b00010000;
	assign font[9][37] = 8'b00010000;
	assign font[10][37] = 8'b00011100;
	assign font[11][37] = 8'b00101100;
	assign font[12][37] = 8'b00101100;
	assign font[13][37] = 8'b00101100;
	assign font[14][37] = 8'b00000000;
	assign font[15][37] = 8'b00000000;

	assign font[0][38] = 8'b00000000;
	assign font[1][38] = 8'b00000000;
	assign font[2][38] = 8'b00000000;
	assign font[3][38] = 8'b00000000;
	assign font[4][38] = 8'b01110000;
	assign font[5][38] = 8'b01001000;
	assign font[6][38] = 8'b01001000;
	assign font[7][38] = 8'b01110100;
	assign font[8][38] = 8'b01110100;
	assign font[9][38] = 8'b01010100;
	assign font[10][38] = 8'b01001000;
	assign font[11][38] = 8'b01011000;
	assign font[12][38] = 8'b01010100;
	assign font[13][38] = 8'b01110100;
	assign font[14][38] = 8'b00000000;
	assign font[15][38] = 8'b00000000;

	assign font[0][39] = 8'b00000000;
	assign font[1][39] = 8'b00000000;
	assign font[2][39] = 8'b00000000;
	assign font[3][39] = 8'b00010000;
	assign font[4][39] = 8'b00100000;
	assign font[5][39] = 8'b00100000;
	assign font[6][39] = 8'b00000000;
	assign font[7][39] = 8'b00000000;
	assign font[8][39] = 8'b00000000;
	assign font[9][39] = 8'b00000000;
	assign font[10][39] = 8'b00000000;
	assign font[11][39] = 8'b00000000;
	assign font[12][39] = 8'b00000000;
	assign font[13][39] = 8'b00000000;
	assign font[14][39] = 8'b00000000;
	assign font[15][39] = 8'b00000000;

	assign font[0][40] = 8'b00000000;
	assign font[1][40] = 8'b00000000;
	assign font[2][40] = 8'b00000000;
	assign font[3][40] = 8'b00000000;
	assign font[4][40] = 8'b00011000;
	assign font[5][40] = 8'b00100000;
	assign font[6][40] = 8'b00100000;
	assign font[7][40] = 8'b00100000;
	assign font[8][40] = 8'b00100000;
	assign font[9][40] = 8'b00100000;
	assign font[10][40] = 8'b00100000;
	assign font[11][40] = 8'b00100000;
	assign font[12][40] = 8'b00100000;
	assign font[13][40] = 8'b00010000;
	assign font[14][40] = 8'b00001000;
	assign font[15][40] = 8'b00000000;

	assign font[0][41] = 8'b00000000;
	assign font[1][41] = 8'b00000000;
	assign font[2][41] = 8'b00000000;
	assign font[3][41] = 8'b00000000;
	assign font[4][41] = 8'b00110000;
	assign font[5][41] = 8'b00010000;
	assign font[6][41] = 8'b00010000;
	assign font[7][41] = 8'b00011000;
	assign font[8][41] = 8'b00011000;
	assign font[9][41] = 8'b00011000;
	assign font[10][41] = 8'b00011000;
	assign font[11][41] = 8'b00010000;
	assign font[12][41] = 8'b00010000;
	assign font[13][41] = 8'b00010000;
	assign font[14][41] = 8'b00100000;
	assign font[15][41] = 8'b00100000;

	assign font[0][42] = 8'b00000000;
	assign font[1][42] = 8'b00000000;
	assign font[2][42] = 8'b00000000;
	assign font[3][42] = 8'b00000000;
	assign font[4][42] = 8'b00000000;
	assign font[5][42] = 8'b00000000;
	assign font[6][42] = 8'b00010000;
	assign font[7][42] = 8'b01011000;
	assign font[8][42] = 8'b00010000;
	assign font[9][42] = 8'b00110000;
	assign font[10][42] = 8'b01011000;
	assign font[11][42] = 8'b00010000;
	assign font[12][42] = 8'b00010000;
	assign font[13][42] = 8'b00000000;
	assign font[14][42] = 8'b00000000;
	assign font[15][42] = 8'b00000000;

	assign font[0][43] = 8'b00000000;
	assign font[1][43] = 8'b00000000;
	assign font[2][43] = 8'b00000000;
	assign font[3][43] = 8'b00000000;
	assign font[4][43] = 8'b00000000;
	assign font[5][43] = 8'b00000000;
	assign font[6][43] = 8'b00011000;
	assign font[7][43] = 8'b00010000;
	assign font[8][43] = 8'b01111100;
	assign font[9][43] = 8'b00010000;
	assign font[10][43] = 8'b00010000;
	assign font[11][43] = 8'b00011000;
	assign font[12][43] = 8'b00000000;
	assign font[13][43] = 8'b00000000;
	assign font[14][43] = 8'b00000000;
	assign font[15][43] = 8'b00000000;

	assign font[0][44] = 8'b00000000;
	assign font[1][44] = 8'b00000000;
	assign font[2][44] = 8'b00000000;
	assign font[3][44] = 8'b00000000;
	assign font[4][44] = 8'b00000000;
	assign font[5][44] = 8'b00000000;
	assign font[6][44] = 8'b00000000;
	assign font[7][44] = 8'b00000000;
	assign font[8][44] = 8'b00000000;
	assign font[9][44] = 8'b00000000;
	assign font[10][44] = 8'b00000000;
	assign font[11][44] = 8'b00000000;
	assign font[12][44] = 8'b00001000;
	assign font[13][44] = 8'b00001000;
	assign font[14][44] = 8'b00011000;
	assign font[15][44] = 8'b00110000;

	assign font[0][45] = 8'b00000000;
	assign font[1][45] = 8'b00000000;
	assign font[2][45] = 8'b00000000;
	assign font[3][45] = 8'b00000000;
	assign font[4][45] = 8'b00000000;
	assign font[5][45] = 8'b00000000;
	assign font[6][45] = 8'b00000000;
	assign font[7][45] = 8'b00000000;
	assign font[8][45] = 8'b00111100;
	assign font[9][45] = 8'b00000000;
	assign font[10][45] = 8'b00000000;
	assign font[11][45] = 8'b00000000;
	assign font[12][45] = 8'b00000000;
	assign font[13][45] = 8'b00000000;
	assign font[14][45] = 8'b00000000;
	assign font[15][45] = 8'b00000000;

	assign font[0][46] = 8'b00000000;
	assign font[1][46] = 8'b00000000;
	assign font[2][46] = 8'b00000000;
	assign font[3][46] = 8'b00000000;
	assign font[4][46] = 8'b00000000;
	assign font[5][46] = 8'b00000000;
	assign font[6][46] = 8'b00000000;
	assign font[7][46] = 8'b00000000;
	assign font[8][46] = 8'b00000000;
	assign font[9][46] = 8'b00000000;
	assign font[10][46] = 8'b00000000;
	assign font[11][46] = 8'b00000000;
	assign font[12][46] = 8'b00011000;
	assign font[13][46] = 8'b00011000;
	assign font[14][46] = 8'b00000000;
	assign font[15][46] = 8'b00000000;

	assign font[0][47] = 8'b00000000;
	assign font[1][47] = 8'b00000000;
	assign font[2][47] = 8'b00000000;
	assign font[3][47] = 8'b00000000;
	assign font[4][47] = 8'b00000100;
	assign font[5][47] = 8'b00000100;
	assign font[6][47] = 8'b00001100;
	assign font[7][47] = 8'b00001000;
	assign font[8][47] = 8'b00001000;
	assign font[9][47] = 8'b00011000;
	assign font[10][47] = 8'b00011000;
	assign font[11][47] = 8'b00110000;
	assign font[12][47] = 8'b00110000;
	assign font[13][47] = 8'b00100000;
	assign font[14][47] = 8'b00100000;
	assign font[15][47] = 8'b00000000;

	assign font[0][48] = 8'b00000000;
	assign font[1][48] = 8'b00000000;
	assign font[2][48] = 8'b00000000;
	assign font[3][48] = 8'b00000000;
	assign font[4][48] = 8'b00110000;
	assign font[5][48] = 8'b00000000;
	assign font[6][48] = 8'b01001000;
	assign font[7][48] = 8'b01001100;
	assign font[8][48] = 8'b01001000;
	assign font[9][48] = 8'b01001000;
	assign font[10][48] = 8'b01001100;
	assign font[11][48] = 8'b01001000;
	assign font[12][48] = 8'b00000000;
	assign font[13][48] = 8'b00110000;
	assign font[14][48] = 8'b00000000;
	assign font[15][48] = 8'b00000000;

	assign font[0][49] = 8'b00000000;
	assign font[1][49] = 8'b00000000;
	assign font[2][49] = 8'b00000000;
	assign font[3][49] = 8'b00000000;
	assign font[4][49] = 8'b00011000;
	assign font[5][49] = 8'b00011000;
	assign font[6][49] = 8'b00011000;
	assign font[7][49] = 8'b00011000;
	assign font[8][49] = 8'b00001000;
	assign font[9][49] = 8'b00001000;
	assign font[10][49] = 8'b00011000;
	assign font[11][49] = 8'b00001000;
	assign font[12][49] = 8'b00001000;
	assign font[13][49] = 8'b00111100;
	assign font[14][49] = 8'b00000000;
	assign font[15][49] = 8'b00000000;

	assign font[0][50] = 8'b00000000;
	assign font[1][50] = 8'b00000000;
	assign font[2][50] = 8'b00000000;
	assign font[3][50] = 8'b00000000;
	assign font[4][50] = 8'b00111000;
	assign font[5][50] = 8'b01001000;
	assign font[6][50] = 8'b01001100;
	assign font[7][50] = 8'b00001100;
	assign font[8][50] = 8'b00011000;
	assign font[9][50] = 8'b00011000;
	assign font[10][50] = 8'b00010000;
	assign font[11][50] = 8'b00100000;
	assign font[12][50] = 8'b00100000;
	assign font[13][50] = 8'b01111000;
	assign font[14][50] = 8'b00000000;
	assign font[15][50] = 8'b00000000;

	assign font[0][51] = 8'b00000000;
	assign font[1][51] = 8'b00000000;
	assign font[2][51] = 8'b00000000;
	assign font[3][51] = 8'b00000000;
	assign font[4][51] = 8'b00111000;
	assign font[5][51] = 8'b01001000;
	assign font[6][51] = 8'b01001100;
	assign font[7][51] = 8'b00001100;
	assign font[8][51] = 8'b00001000;
	assign font[9][51] = 8'b00111000;
	assign font[10][51] = 8'b00001100;
	assign font[11][51] = 8'b00001100;
	assign font[12][51] = 8'b00001000;
	assign font[13][51] = 8'b00111000;
	assign font[14][51] = 8'b00000000;
	assign font[15][51] = 8'b00000000;

	assign font[0][52] = 8'b00000000;
	assign font[1][52] = 8'b00000000;
	assign font[2][52] = 8'b00000000;
	assign font[3][52] = 8'b00000000;
	assign font[4][52] = 8'b00011000;
	assign font[5][52] = 8'b00001000;
	assign font[6][52] = 8'b00101000;
	assign font[7][52] = 8'b00101000;
	assign font[8][52] = 8'b00101000;
	assign font[9][52] = 8'b01001100;
	assign font[10][52] = 8'b01111100;
	assign font[11][52] = 8'b00001000;
	assign font[12][52] = 8'b00001000;
	assign font[13][52] = 8'b00001100;
	assign font[14][52] = 8'b00000000;
	assign font[15][52] = 8'b00000000;

	assign font[0][53] = 8'b00000000;
	assign font[1][53] = 8'b00000000;
	assign font[2][53] = 8'b00000000;
	assign font[3][53] = 8'b00000000;
	assign font[4][53] = 8'b01111100;
	assign font[5][53] = 8'b01100000;
	assign font[6][53] = 8'b01100000;
	assign font[7][53] = 8'b01111000;
	assign font[8][53] = 8'b01101000;
	assign font[9][53] = 8'b01101100;
	assign font[10][53] = 8'b00000100;
	assign font[11][53] = 8'b00000100;
	assign font[12][53] = 8'b01001100;
	assign font[13][53] = 8'b00111000;
	assign font[14][53] = 8'b00000000;
	assign font[15][53] = 8'b00000000;

	assign font[0][54] = 8'b00000000;
	assign font[1][54] = 8'b00000000;
	assign font[2][54] = 8'b00000000;
	assign font[3][54] = 8'b00000000;
	assign font[4][54] = 8'b00011000;
	assign font[5][54] = 8'b00000000;
	assign font[6][54] = 8'b00100000;
	assign font[7][54] = 8'b01100000;
	assign font[8][54] = 8'b00100000;
	assign font[9][54] = 8'b00111100;
	assign font[10][54] = 8'b00100110;
	assign font[11][54] = 8'b00100100;
	assign font[12][54] = 8'b00000100;
	assign font[13][54] = 8'b00011100;
	assign font[14][54] = 8'b00000000;
	assign font[15][54] = 8'b00000000;

	assign font[0][55] = 8'b00000000;
	assign font[1][55] = 8'b00000000;
	assign font[2][55] = 8'b00000000;
	assign font[3][55] = 8'b00000000;
	assign font[4][55] = 8'b01111100;
	assign font[5][55] = 8'b00001000;
	assign font[6][55] = 8'b00001000;
	assign font[7][55] = 8'b00001000;
	assign font[8][55] = 8'b00010000;
	assign font[9][55] = 8'b00011000;
	assign font[10][55] = 8'b00011000;
	assign font[11][55] = 8'b00010000;
	assign font[12][55] = 8'b00110000;
	assign font[13][55] = 8'b00100000;
	assign font[14][55] = 8'b00000000;
	assign font[15][55] = 8'b00000000;

	assign font[0][56] = 8'b00000000;
	assign font[1][56] = 8'b00000000;
	assign font[2][56] = 8'b00000000;
	assign font[3][56] = 8'b00000000;
	assign font[4][56] = 8'b00111000;
	assign font[5][56] = 8'b01001000;
	assign font[6][56] = 8'b01001100;
	assign font[7][56] = 8'b01001000;
	assign font[8][56] = 8'b01001000;
	assign font[9][56] = 8'b00111000;
	assign font[10][56] = 8'b01001100;
	assign font[11][56] = 8'b01001000;
	assign font[12][56] = 8'b01001000;
	assign font[13][56] = 8'b00111000;
	assign font[14][56] = 8'b00000000;
	assign font[15][56] = 8'b00000000;

	assign font[0][57] = 8'b00000000;
	assign font[1][57] = 8'b00000000;
	assign font[2][57] = 8'b00000000;
	assign font[3][57] = 8'b00000000;
	assign font[4][57] = 8'b00111000;
	assign font[5][57] = 8'b01001000;
	assign font[6][57] = 8'b01000100;
	assign font[7][57] = 8'b01000100;
	assign font[8][57] = 8'b01000100;
	assign font[9][57] = 8'b00111100;
	assign font[10][57] = 8'b00000100;
	assign font[11][57] = 8'b00001000;
	assign font[12][57] = 8'b00001000;
	assign font[13][57] = 8'b00111000;
	assign font[14][57] = 8'b00000000;
	assign font[15][57] = 8'b00000000;

	assign font[0][58] = 8'b00000000;
	assign font[1][58] = 8'b00000000;
	assign font[2][58] = 8'b00000000;
	assign font[3][58] = 8'b00000000;
	assign font[4][58] = 8'b00000000;
	assign font[5][58] = 8'b00000000;
	assign font[6][58] = 8'b00000000;
	assign font[7][58] = 8'b00011000;
	assign font[8][58] = 8'b00011000;
	assign font[9][58] = 8'b00000000;
	assign font[10][58] = 8'b00000000;
	assign font[11][58] = 8'b00000000;
	assign font[12][58] = 8'b00011000;
	assign font[13][58] = 8'b00011000;
	assign font[14][58] = 8'b00000000;
	assign font[15][58] = 8'b00000000;

	assign font[0][59] = 8'b00000000;
	assign font[1][59] = 8'b00000000;
	assign font[2][59] = 8'b00000000;
	assign font[3][59] = 8'b00000000;
	assign font[4][59] = 8'b00000000;
	assign font[5][59] = 8'b00000000;
	assign font[6][59] = 8'b00010000;
	assign font[7][59] = 8'b00010000;
	assign font[8][59] = 8'b00000000;
	assign font[9][59] = 8'b00000000;
	assign font[10][59] = 8'b00000000;
	assign font[11][59] = 8'b00010000;
	assign font[12][59] = 8'b00010000;
	assign font[13][59] = 8'b00011000;
	assign font[14][59] = 8'b00110000;
	assign font[15][59] = 8'b01100000;

	assign font[0][60] = 8'b00000000;
	assign font[1][60] = 8'b00000000;
	assign font[2][60] = 8'b00000000;
	assign font[3][60] = 8'b00000000;
	assign font[4][60] = 8'b00001100;
	assign font[5][60] = 8'b00001000;
	assign font[6][60] = 8'b00001000;
	assign font[7][60] = 8'b00010000;
	assign font[8][60] = 8'b00100000;
	assign font[9][60] = 8'b00100000;
	assign font[10][60] = 8'b00010000;
	assign font[11][60] = 8'b00001000;
	assign font[12][60] = 8'b00001000;
	assign font[13][60] = 8'b00001100;
	assign font[14][60] = 8'b00000000;
	assign font[15][60] = 8'b00000000;

	assign font[0][61] = 8'b00000000;
	assign font[1][61] = 8'b00000000;
	assign font[2][61] = 8'b00000000;
	assign font[3][61] = 8'b00000000;
	assign font[4][61] = 8'b00000000;
	assign font[5][61] = 8'b00000000;
	assign font[6][61] = 8'b00000000;
	assign font[7][61] = 8'b00111100;
	assign font[8][61] = 8'b00000000;
	assign font[9][61] = 8'b00000000;
	assign font[10][61] = 8'b00111100;
	assign font[11][61] = 8'b00000000;
	assign font[12][61] = 8'b00000000;
	assign font[13][61] = 8'b00000000;
	assign font[14][61] = 8'b00000000;
	assign font[15][61] = 8'b00000000;

	assign font[0][62] = 8'b00000000;
	assign font[1][62] = 8'b00000000;
	assign font[2][62] = 8'b00000000;
	assign font[3][62] = 8'b00000000;
	assign font[4][62] = 8'b01000000;
	assign font[5][62] = 8'b01000000;
	assign font[6][62] = 8'b00100000;
	assign font[7][62] = 8'b00010000;
	assign font[8][62] = 8'b00010000;
	assign font[9][62] = 8'b00011000;
	assign font[10][62] = 8'b00010000;
	assign font[11][62] = 8'b00100000;
	assign font[12][62] = 8'b00100000;
	assign font[13][62] = 8'b01000000;
	assign font[14][62] = 8'b00000000;
	assign font[15][62] = 8'b00000000;

	assign font[0][63] = 8'b00000000;
	assign font[1][63] = 8'b00000000;
	assign font[2][63] = 8'b00000000;
	assign font[3][63] = 8'b00000000;
	assign font[4][63] = 8'b00111000;
	assign font[5][63] = 8'b00101000;
	assign font[6][63] = 8'b01101000;
	assign font[7][63] = 8'b00001000;
	assign font[8][63] = 8'b00011000;
	assign font[9][63] = 8'b00010000;
	assign font[10][63] = 8'b00010000;
	assign font[11][63] = 8'b00000000;
	assign font[12][63] = 8'b00000000;
	assign font[13][63] = 8'b00010000;
	assign font[14][63] = 8'b00000000;
	assign font[15][63] = 8'b00000000;

	assign font[0][64] = 8'b00000000;
	assign font[1][64] = 8'b00000000;
	assign font[2][64] = 8'b00000000;
	assign font[3][64] = 8'b00000000;
	assign font[4][64] = 8'b00111100;
	assign font[5][64] = 8'b00101100;
	assign font[6][64] = 8'b01011110;
	assign font[7][64] = 8'b01010100;
	assign font[8][64] = 8'b01010100;
	assign font[9][64] = 8'b01010110;
	assign font[10][64] = 8'b01011100;
	assign font[11][64] = 8'b00100000;
	assign font[12][64] = 8'b00100000;
	assign font[13][64] = 8'b00111100;
	assign font[14][64] = 8'b00000000;
	assign font[15][64] = 8'b00000000;

	assign font[0][65] = 8'b00000000;
	assign font[1][65] = 8'b00000000;
	assign font[2][65] = 8'b00000000;
	assign font[3][65] = 8'b00000000;
	assign font[4][65] = 8'b00110000;
	assign font[5][65] = 8'b00111000;
	assign font[6][65] = 8'b00101000;
	assign font[7][65] = 8'b01101000;
	assign font[8][65] = 8'b01001000;
	assign font[9][65] = 8'b01101000;
	assign font[10][65] = 8'b01111000;
	assign font[11][65] = 8'b01001000;
	assign font[12][65] = 8'b01000100;
	assign font[13][65] = 8'b01000100;
	assign font[14][65] = 8'b00000000;
	assign font[15][65] = 8'b00000000;

	assign font[0][66] = 8'b00000000;
	assign font[1][66] = 8'b00000000;
	assign font[2][66] = 8'b00000000;
	assign font[3][66] = 8'b00000000;
	assign font[4][66] = 8'b01111100;
	assign font[5][66] = 8'b01000100;
	assign font[6][66] = 8'b01000100;
	assign font[7][66] = 8'b01000100;
	assign font[8][66] = 8'b01000100;
	assign font[9][66] = 8'b01111100;
	assign font[10][66] = 8'b01000100;
	assign font[11][66] = 8'b01000100;
	assign font[12][66] = 8'b01100100;
	assign font[13][66] = 8'b01111100;
	assign font[14][66] = 8'b00000000;
	assign font[15][66] = 8'b00000000;

	assign font[0][67] = 8'b00000000;
	assign font[1][67] = 8'b00000000;
	assign font[2][67] = 8'b00000000;
	assign font[3][67] = 8'b00000000;
	assign font[4][67] = 8'b00111000;
	assign font[5][67] = 8'b00101000;
	assign font[6][67] = 8'b00100100;
	assign font[7][67] = 8'b01000000;
	assign font[8][67] = 8'b01000000;
	assign font[9][67] = 8'b01000000;
	assign font[10][67] = 8'b01000000;
	assign font[11][67] = 8'b01000000;
	assign font[12][67] = 8'b01000100;
	assign font[13][67] = 8'b00111000;
	assign font[14][67] = 8'b00000000;
	assign font[15][67] = 8'b00000000;

	assign font[0][68] = 8'b00000000;
	assign font[1][68] = 8'b00000000;
	assign font[2][68] = 8'b00000000;
	assign font[3][68] = 8'b00000000;
	assign font[4][68] = 8'b01111000;
	assign font[5][68] = 8'b01001000;
	assign font[6][68] = 8'b01001100;
	assign font[7][68] = 8'b01000110;
	assign font[8][68] = 8'b01000100;
	assign font[9][68] = 8'b01100100;
	assign font[10][68] = 8'b01000110;
	assign font[11][68] = 8'b01001100;
	assign font[12][68] = 8'b01101000;
	assign font[13][68] = 8'b01111000;
	assign font[14][68] = 8'b00000000;
	assign font[15][68] = 8'b00000000;

	assign font[0][69] = 8'b00000000;
	assign font[1][69] = 8'b00000000;
	assign font[2][69] = 8'b00000000;
	assign font[3][69] = 8'b00000000;
	assign font[4][69] = 8'b00111100;
	assign font[5][69] = 8'b00100000;
	assign font[6][69] = 8'b00100000;
	assign font[7][69] = 8'b00100000;
	assign font[8][69] = 8'b00100000;
	assign font[9][69] = 8'b00111100;
	assign font[10][69] = 8'b00100000;
	assign font[11][69] = 8'b00100000;
	assign font[12][69] = 8'b00110000;
	assign font[13][69] = 8'b00111100;
	assign font[14][69] = 8'b00000000;
	assign font[15][69] = 8'b00000000;

	assign font[0][70] = 8'b00000000;
	assign font[1][70] = 8'b00000000;
	assign font[2][70] = 8'b00000000;
	assign font[3][70] = 8'b00000000;
	assign font[4][70] = 8'b00111100;
	assign font[5][70] = 8'b00100000;
	assign font[6][70] = 8'b00100000;
	assign font[7][70] = 8'b00100000;
	assign font[8][70] = 8'b00100000;
	assign font[9][70] = 8'b00111100;
	assign font[10][70] = 8'b00100000;
	assign font[11][70] = 8'b00100000;
	assign font[12][70] = 8'b00100000;
	assign font[13][70] = 8'b00110000;
	assign font[14][70] = 8'b00000000;
	assign font[15][70] = 8'b00000000;

	assign font[0][71] = 8'b00000000;
	assign font[1][71] = 8'b00000000;
	assign font[2][71] = 8'b00000000;
	assign font[3][71] = 8'b00000000;
	assign font[4][71] = 8'b00111000;
	assign font[5][71] = 8'b00101000;
	assign font[6][71] = 8'b00100100;
	assign font[7][71] = 8'b01000000;
	assign font[8][71] = 8'b01000000;
	assign font[9][71] = 8'b01001100;
	assign font[10][71] = 8'b01000100;
	assign font[11][71] = 8'b01000100;
	assign font[12][71] = 8'b01000110;
	assign font[13][71] = 8'b00111000;
	assign font[14][71] = 8'b00000000;
	assign font[15][71] = 8'b00000000;

	assign font[0][72] = 8'b00000000;
	assign font[1][72] = 8'b00000000;
	assign font[2][72] = 8'b00000000;
	assign font[3][72] = 8'b00000000;
	assign font[4][72] = 8'b01100110;
	assign font[5][72] = 8'b01000100;
	assign font[6][72] = 8'b01100110;
	assign font[7][72] = 8'b01000100;
	assign font[8][72] = 8'b01100110;
	assign font[9][72] = 8'b01111100;
	assign font[10][72] = 8'b01000100;
	assign font[11][72] = 8'b01000100;
	assign font[12][72] = 8'b01000110;
	assign font[13][72] = 8'b01100110;
	assign font[14][72] = 8'b00000000;
	assign font[15][72] = 8'b00000000;

	assign font[0][73] = 8'b00000000;
	assign font[1][73] = 8'b00000000;
	assign font[2][73] = 8'b00000000;
	assign font[3][73] = 8'b00000000;
	assign font[4][73] = 8'b00111000;
	assign font[5][73] = 8'b00011000;
	assign font[6][73] = 8'b00010000;
	assign font[7][73] = 8'b00010000;
	assign font[8][73] = 8'b00010000;
	assign font[9][73] = 8'b00011000;
	assign font[10][73] = 8'b00010000;
	assign font[11][73] = 8'b00010000;
	assign font[12][73] = 8'b00011000;
	assign font[13][73] = 8'b00111000;
	assign font[14][73] = 8'b00000000;
	assign font[15][73] = 8'b00000000;

	assign font[0][74] = 8'b00000000;
	assign font[1][74] = 8'b00000000;
	assign font[2][74] = 8'b00000000;
	assign font[3][74] = 8'b00000000;
	assign font[4][74] = 8'b00011100;
	assign font[5][74] = 8'b00001000;
	assign font[6][74] = 8'b00001000;
	assign font[7][74] = 8'b00001000;
	assign font[8][74] = 8'b00001000;
	assign font[9][74] = 8'b00001100;
	assign font[10][74] = 8'b00001000;
	assign font[11][74] = 8'b01001000;
	assign font[12][74] = 8'b01101100;
	assign font[13][74] = 8'b00111000;
	assign font[14][74] = 8'b00000000;
	assign font[15][74] = 8'b00000000;

	assign font[0][75] = 8'b00000000;
	assign font[1][75] = 8'b00000000;
	assign font[2][75] = 8'b00000000;
	assign font[3][75] = 8'b00000000;
	assign font[4][75] = 8'b01001000;
	assign font[5][75] = 8'b01001000;
	assign font[6][75] = 8'b01010000;
	assign font[7][75] = 8'b01010000;
	assign font[8][75] = 8'b01100000;
	assign font[9][75] = 8'b01100000;
	assign font[10][75] = 8'b01010000;
	assign font[11][75] = 8'b01010000;
	assign font[12][75] = 8'b01001000;
	assign font[13][75] = 8'b01001000;
	assign font[14][75] = 8'b00000000;
	assign font[15][75] = 8'b00000000;

	assign font[0][76] = 8'b00000000;
	assign font[1][76] = 8'b00000000;
	assign font[2][76] = 8'b00000000;
	assign font[3][76] = 8'b00000000;
	assign font[4][76] = 8'b01000000;
	assign font[5][76] = 8'b01000000;
	assign font[6][76] = 8'b01000000;
	assign font[7][76] = 8'b01000000;
	assign font[8][76] = 8'b01000000;
	assign font[9][76] = 8'b01100000;
	assign font[10][76] = 8'b01000000;
	assign font[11][76] = 8'b01000000;
	assign font[12][76] = 8'b01100000;
	assign font[13][76] = 8'b01111100;
	assign font[14][76] = 8'b00000000;
	assign font[15][76] = 8'b00000000;

	assign font[0][77] = 8'b00000000;
	assign font[1][77] = 8'b00000000;
	assign font[2][77] = 8'b00000000;
	assign font[3][77] = 8'b00000000;
	assign font[4][77] = 8'b01101100;
	assign font[5][77] = 8'b01101100;
	assign font[6][77] = 8'b01110100;
	assign font[7][77] = 8'b01101100;
	assign font[8][77] = 8'b01101100;
	assign font[9][77] = 8'b01011100;
	assign font[10][77] = 8'b01010110;
	assign font[11][77] = 8'b01010100;
	assign font[12][77] = 8'b01111100;
	assign font[13][77] = 8'b01100110;
	assign font[14][77] = 8'b00000000;
	assign font[15][77] = 8'b00000000;

	assign font[0][78] = 8'b00000000;
	assign font[1][78] = 8'b00000000;
	assign font[2][78] = 8'b00000000;
	assign font[3][78] = 8'b00000000;
	assign font[4][78] = 8'b01000100;
	assign font[5][78] = 8'b01100100;
	assign font[6][78] = 8'b01100100;
	assign font[7][78] = 8'b01110100;
	assign font[8][78] = 8'b01010100;
	assign font[9][78] = 8'b01010100;
	assign font[10][78] = 8'b01001100;
	assign font[11][78] = 8'b01001100;
	assign font[12][78] = 8'b01000100;
	assign font[13][78] = 8'b01000100;
	assign font[14][78] = 8'b00000000;
	assign font[15][78] = 8'b00000000;

	assign font[0][79] = 8'b00000000;
	assign font[1][79] = 8'b00000000;
	assign font[2][79] = 8'b00000000;
	assign font[3][79] = 8'b00000000;
	assign font[4][79] = 8'b00111000;
	assign font[5][79] = 8'b00101000;
	assign font[6][79] = 8'b00101100;
	assign font[7][79] = 8'b01000110;
	assign font[8][79] = 8'b01000100;
	assign font[9][79] = 8'b01000100;
	assign font[10][79] = 8'b01000110;
	assign font[11][79] = 8'b00101100;
	assign font[12][79] = 8'b00101000;
	assign font[13][79] = 8'b00111000;
	assign font[14][79] = 8'b00000000;
	assign font[15][79] = 8'b00000000;

	assign font[0][80] = 8'b00000000;
	assign font[1][80] = 8'b00000000;
	assign font[2][80] = 8'b00000000;
	assign font[3][80] = 8'b00000000;
	assign font[4][80] = 8'b01111000;
	assign font[5][80] = 8'b01001000;
	assign font[6][80] = 8'b01001100;
	assign font[7][80] = 8'b01001100;
	assign font[8][80] = 8'b01001000;
	assign font[9][80] = 8'b01111000;
	assign font[10][80] = 8'b01000000;
	assign font[11][80] = 8'b01000000;
	assign font[12][80] = 8'b01000000;
	assign font[13][80] = 8'b01100000;
	assign font[14][80] = 8'b00000000;
	assign font[15][80] = 8'b00000000;

	assign font[0][81] = 8'b00000000;
	assign font[1][81] = 8'b00000000;
	assign font[2][81] = 8'b00000000;
	assign font[3][81] = 8'b00000000;
	assign font[4][81] = 8'b00111000;
	assign font[5][81] = 8'b00101000;
	assign font[6][81] = 8'b00101100;
	assign font[7][81] = 8'b01000110;
	assign font[8][81] = 8'b01000100;
	assign font[9][81] = 8'b01000100;
	assign font[10][81] = 8'b01011110;
	assign font[11][81] = 8'b00101100;
	assign font[12][81] = 8'b00101000;
	assign font[13][81] = 8'b00111000;
	assign font[14][81] = 8'b00001100;
	assign font[15][81] = 8'b00000100;

	assign font[0][82] = 8'b00000000;
	assign font[1][82] = 8'b00000000;
	assign font[2][82] = 8'b00000000;
	assign font[3][82] = 8'b00000000;
	assign font[4][82] = 8'b01111100;
	assign font[5][82] = 8'b01001100;
	assign font[6][82] = 8'b01001100;
	assign font[7][82] = 8'b01001100;
	assign font[8][82] = 8'b01001100;
	assign font[9][82] = 8'b01111000;
	assign font[10][82] = 8'b01101100;
	assign font[11][82] = 8'b01001100;
	assign font[12][82] = 8'b01001100;
	assign font[13][82] = 8'b01100100;
	assign font[14][82] = 8'b00000000;
	assign font[15][82] = 8'b00000000;

	assign font[0][83] = 8'b00000000;
	assign font[1][83] = 8'b00000000;
	assign font[2][83] = 8'b00000000;
	assign font[3][83] = 8'b00000000;
	assign font[4][83] = 8'b00111000;
	assign font[5][83] = 8'b01001000;
	assign font[6][83] = 8'b01001100;
	assign font[7][83] = 8'b01000000;
	assign font[8][83] = 8'b01000000;
	assign font[9][83] = 8'b00111000;
	assign font[10][83] = 8'b00001100;
	assign font[11][83] = 8'b00001100;
	assign font[12][83] = 8'b00001000;
	assign font[13][83] = 8'b00111000;
	assign font[14][83] = 8'b00000000;
	assign font[15][83] = 8'b00000000;

	assign font[0][84] = 8'b00000000;
	assign font[1][84] = 8'b00000000;
	assign font[2][84] = 8'b00000000;
	assign font[3][84] = 8'b00000000;
	assign font[4][84] = 8'b01111100;
	assign font[5][84] = 8'b00010000;
	assign font[6][84] = 8'b00010000;
	assign font[7][84] = 8'b00011000;
	assign font[8][84] = 8'b00010000;
	assign font[9][84] = 8'b00010000;
	assign font[10][84] = 8'b00011000;
	assign font[11][84] = 8'b00010000;
	assign font[12][84] = 8'b00010000;
	assign font[13][84] = 8'b00011000;
	assign font[14][84] = 8'b00000000;
	assign font[15][84] = 8'b00000000;

	assign font[0][85] = 8'b00000000;
	assign font[1][85] = 8'b00000000;
	assign font[2][85] = 8'b00000000;
	assign font[3][85] = 8'b00000000;
	assign font[4][85] = 8'b01100100;
	assign font[5][85] = 8'b01000100;
	assign font[6][85] = 8'b01100100;
	assign font[7][85] = 8'b01001100;
	assign font[8][85] = 8'b01000100;
	assign font[9][85] = 8'b01000100;
	assign font[10][85] = 8'b01001110;
	assign font[11][85] = 8'b01000110;
	assign font[12][85] = 8'b01001000;
	assign font[13][85] = 8'b00111000;
	assign font[14][85] = 8'b00000000;
	assign font[15][85] = 8'b00000000;

	assign font[0][86] = 8'b00000000;
	assign font[1][86] = 8'b00000000;
	assign font[2][86] = 8'b00000000;
	assign font[3][86] = 8'b00000000;
	assign font[4][86] = 8'b01101100;
	assign font[5][86] = 8'b01001100;
	assign font[6][86] = 8'b01001100;
	assign font[7][86] = 8'b01101100;
	assign font[8][86] = 8'b00101000;
	assign font[9][86] = 8'b00101000;
	assign font[10][86] = 8'b00101000;
	assign font[11][86] = 8'b00111000;
	assign font[12][86] = 8'b00111000;
	assign font[13][86] = 8'b00010000;
	assign font[14][86] = 8'b00000000;
	assign font[15][86] = 8'b00000000;

	assign font[0][87] = 8'b00000000;
	assign font[1][87] = 8'b00000000;
	assign font[2][87] = 8'b00000000;
	assign font[3][87] = 8'b00000000;
	assign font[4][87] = 8'b01110110;
	assign font[5][87] = 8'b01010100;
	assign font[6][87] = 8'b01010100;
	assign font[7][87] = 8'b01010100;
	assign font[8][87] = 8'b01010110;
	assign font[9][87] = 8'b01010100;
	assign font[10][87] = 8'b01011100;
	assign font[11][87] = 8'b01011100;
	assign font[12][87] = 8'b00101000;
	assign font[13][87] = 8'b00101000;
	assign font[14][87] = 8'b00000000;
	assign font[15][87] = 8'b00000000;

	assign font[0][88] = 8'b00000000;
	assign font[1][88] = 8'b00000000;
	assign font[2][88] = 8'b00000000;
	assign font[3][88] = 8'b00000000;
	assign font[4][88] = 8'b01000100;
	assign font[5][88] = 8'b01001100;
	assign font[6][88] = 8'b01001000;
	assign font[7][88] = 8'b00101000;
	assign font[8][88] = 8'b00101000;
	assign font[9][88] = 8'b00110000;
	assign font[10][88] = 8'b00101000;
	assign font[11][88] = 8'b01001000;
	assign font[12][88] = 8'b01001100;
	assign font[13][88] = 8'b11001100;
	assign font[14][88] = 8'b00000000;
	assign font[15][88] = 8'b00000000;

	assign font[0][89] = 8'b00000000;
	assign font[1][89] = 8'b00000000;
	assign font[2][89] = 8'b00000000;
	assign font[3][89] = 8'b00000000;
	assign font[4][89] = 8'b01001100;
	assign font[5][89] = 8'b01001100;
	assign font[6][89] = 8'b01001000;
	assign font[7][89] = 8'b01001100;
	assign font[8][89] = 8'b01101000;
	assign font[9][89] = 8'b00110000;
	assign font[10][89] = 8'b00110000;
	assign font[11][89] = 8'b00110000;
	assign font[12][89] = 8'b00110000;
	assign font[13][89] = 8'b00110000;
	assign font[14][89] = 8'b00000000;
	assign font[15][89] = 8'b00000000;

	assign font[0][90] = 8'b00000000;
	assign font[1][90] = 8'b00000000;
	assign font[2][90] = 8'b00000000;
	assign font[3][90] = 8'b00000000;
	assign font[4][90] = 8'b01111100;
	assign font[5][90] = 8'b00001000;
	assign font[6][90] = 8'b00001000;
	assign font[7][90] = 8'b00011000;
	assign font[8][90] = 8'b00011000;
	assign font[9][90] = 8'b00010000;
	assign font[10][90] = 8'b00100000;
	assign font[11][90] = 8'b00100000;
	assign font[12][90] = 8'b01000000;
	assign font[13][90] = 8'b01111000;
	assign font[14][90] = 8'b00000000;
	assign font[15][90] = 8'b00000000;

	assign font[0][91] = 8'b00000000;
	assign font[1][91] = 8'b00000000;
	assign font[2][91] = 8'b00000000;
	assign font[3][91] = 8'b00011000;
	assign font[4][91] = 8'b00011000;
	assign font[5][91] = 8'b00010000;
	assign font[6][91] = 8'b00011000;
	assign font[7][91] = 8'b00010000;
	assign font[8][91] = 8'b00010000;
	assign font[9][91] = 8'b00010000;
	assign font[10][91] = 8'b00011000;
	assign font[11][91] = 8'b00010000;
	assign font[12][91] = 8'b00010000;
	assign font[13][91] = 8'b00011000;
	assign font[14][91] = 8'b00011000;
	assign font[15][91] = 8'b00000000;

	assign font[0][92] = 8'b00000000;
	assign font[1][92] = 8'b00000000;
	assign font[2][92] = 8'b00000000;
	assign font[3][92] = 8'b00000000;
	assign font[4][92] = 8'b01100000;
	assign font[5][92] = 8'b00100000;
	assign font[6][92] = 8'b00100000;
	assign font[7][92] = 8'b00110000;
	assign font[8][92] = 8'b00010000;
	assign font[9][92] = 8'b00010000;
	assign font[10][92] = 8'b00011000;
	assign font[11][92] = 8'b00001000;
	assign font[12][92] = 8'b00001000;
	assign font[13][92] = 8'b00001100;
	assign font[14][92] = 8'b00001100;
	assign font[15][92] = 8'b00000000;

	assign font[0][93] = 8'b00000000;
	assign font[1][93] = 8'b00000000;
	assign font[2][93] = 8'b00000000;
	assign font[3][93] = 8'b00011100;
	assign font[4][93] = 8'b00001100;
	assign font[5][93] = 8'b00001100;
	assign font[6][93] = 8'b00001100;
	assign font[7][93] = 8'b00001100;
	assign font[8][93] = 8'b00001100;
	assign font[9][93] = 8'b00001100;
	assign font[10][93] = 8'b00001100;
	assign font[11][93] = 8'b00001100;
	assign font[12][93] = 8'b00001100;
	assign font[13][93] = 8'b00001100;
	assign font[14][93] = 8'b00011100;
	assign font[15][93] = 8'b00000000;

	assign font[0][94] = 8'b00000000;
	assign font[1][94] = 8'b00000000;
	assign font[2][94] = 8'b00000000;
	assign font[3][94] = 8'b00000000;
	assign font[4][94] = 8'b00000000;
	assign font[5][94] = 8'b00011000;
	assign font[6][94] = 8'b00011100;
	assign font[7][94] = 8'b00100100;
	assign font[8][94] = 8'b00100100;
	assign font[9][94] = 8'b00000000;
	assign font[10][94] = 8'b00000000;
	assign font[11][94] = 8'b00000000;
	assign font[12][94] = 8'b00000000;
	assign font[13][94] = 8'b00000000;
	assign font[14][94] = 8'b00000000;
	assign font[15][94] = 8'b00000000;

	assign font[0][95] = 8'b00000000;
	assign font[1][95] = 8'b00000000;
	assign font[2][95] = 8'b00000000;
	assign font[3][95] = 8'b00000000;
	assign font[4][95] = 8'b00000000;
	assign font[5][95] = 8'b00000000;
	assign font[6][95] = 8'b00000000;
	assign font[7][95] = 8'b00000000;
	assign font[8][95] = 8'b00000000;
	assign font[9][95] = 8'b00000000;
	assign font[10][95] = 8'b00000000;
	assign font[11][95] = 8'b00000000;
	assign font[12][95] = 8'b01111100;
	assign font[13][95] = 8'b00000000;
	assign font[14][95] = 8'b00000000;
	assign font[15][95] = 8'b00000000;

	assign font[0][96] = 8'b00000000;
	assign font[1][96] = 8'b00000000;
	assign font[2][96] = 8'b00000000;
	assign font[3][96] = 8'b00000000;
	assign font[4][96] = 8'b00110000;
	assign font[5][96] = 8'b00010000;
	assign font[6][96] = 8'b00000000;
	assign font[7][96] = 8'b00000000;
	assign font[8][96] = 8'b00000000;
	assign font[9][96] = 8'b00000000;
	assign font[10][96] = 8'b00000000;
	assign font[11][96] = 8'b00000000;
	assign font[12][96] = 8'b00000000;
	assign font[13][96] = 8'b00000000;
	assign font[14][96] = 8'b00000000;
	assign font[15][96] = 8'b00000000;

	assign font[0][97] = 8'b00000000;
	assign font[1][97] = 8'b00000000;
	assign font[2][97] = 8'b00000000;
	assign font[3][97] = 8'b00000000;
	assign font[4][97] = 8'b00000000;
	assign font[5][97] = 8'b00000000;
	assign font[6][97] = 8'b00000000;
	assign font[7][97] = 8'b00111000;
	assign font[8][97] = 8'b00001000;
	assign font[9][97] = 8'b00000100;
	assign font[10][97] = 8'b00111100;
	assign font[11][97] = 8'b00100100;
	assign font[12][97] = 8'b00100100;
	assign font[13][97] = 8'b00111110;
	assign font[14][97] = 8'b00000000;
	assign font[15][97] = 8'b00000000;

	assign font[0][98] = 8'b00000000;
	assign font[1][98] = 8'b00000000;
	assign font[2][98] = 8'b00000000;
	assign font[3][98] = 8'b00000000;
	assign font[4][98] = 8'b11000000;
	assign font[5][98] = 8'b01000000;
	assign font[6][98] = 8'b01000000;
	assign font[7][98] = 8'b11011000;
	assign font[8][98] = 8'b11101000;
	assign font[9][98] = 8'b01100100;
	assign font[10][98] = 8'b01000100;
	assign font[11][98] = 8'b11000100;
	assign font[12][98] = 8'b01000000;
	assign font[13][98] = 8'b01111000;
	assign font[14][98] = 8'b00000000;
	assign font[15][98] = 8'b00000000;

	assign font[0][99] = 8'b00000000;
	assign font[1][99] = 8'b00000000;
	assign font[2][99] = 8'b00000000;
	assign font[3][99] = 8'b00000000;
	assign font[4][99] = 8'b00000000;
	assign font[5][99] = 8'b00000000;
	assign font[6][99] = 8'b00000000;
	assign font[7][99] = 8'b00111000;
	assign font[8][99] = 8'b01001000;
	assign font[9][99] = 8'b01001100;
	assign font[10][99] = 8'b01000000;
	assign font[11][99] = 8'b01000000;
	assign font[12][99] = 8'b01001100;
	assign font[13][99] = 8'b00111000;
	assign font[14][99] = 8'b00000000;
	assign font[15][99] = 8'b00000000;

	assign font[0][100] = 8'b00000000;
	assign font[1][100] = 8'b00000000;
	assign font[2][100] = 8'b00000000;
	assign font[3][100] = 8'b00000000;
	assign font[4][100] = 8'b00001100;
	assign font[5][100] = 8'b00000100;
	assign font[6][100] = 8'b00000100;
	assign font[7][100] = 8'b00110100;
	assign font[8][100] = 8'b01000100;
	assign font[9][100] = 8'b01000100;
	assign font[10][100] = 8'b01000100;
	assign font[11][100] = 8'b01000100;
	assign font[12][100] = 8'b01000100;
	assign font[13][100] = 8'b00111100;
	assign font[14][100] = 8'b00000000;
	assign font[15][100] = 8'b00000000;

	assign font[0][101] = 8'b00000000;
	assign font[1][101] = 8'b00000000;
	assign font[2][101] = 8'b00000000;
	assign font[3][101] = 8'b00000000;
	assign font[4][101] = 8'b00000000;
	assign font[5][101] = 8'b00000000;
	assign font[6][101] = 8'b00000000;
	assign font[7][101] = 8'b00111000;
	assign font[8][101] = 8'b01001100;
	assign font[9][101] = 8'b01001100;
	assign font[10][101] = 8'b01111100;
	assign font[11][101] = 8'b01000000;
	assign font[12][101] = 8'b01000000;
	assign font[13][101] = 8'b00111000;
	assign font[14][101] = 8'b00000000;
	assign font[15][101] = 8'b00000000;

	assign font[0][102] = 8'b00000000;
	assign font[1][102] = 8'b00000000;
	assign font[2][102] = 8'b00000000;
	assign font[3][102] = 8'b00000000;
	assign font[4][102] = 8'b00111100;
	assign font[5][102] = 8'b00100000;
	assign font[6][102] = 8'b00100000;
	assign font[7][102] = 8'b01111100;
	assign font[8][102] = 8'b00100000;
	assign font[9][102] = 8'b00100000;
	assign font[10][102] = 8'b00100000;
	assign font[11][102] = 8'b00100000;
	assign font[12][102] = 8'b00110000;
	assign font[13][102] = 8'b01110000;
	assign font[14][102] = 8'b00000000;
	assign font[15][102] = 8'b00000000;

	assign font[0][103] = 8'b00000000;
	assign font[1][103] = 8'b00000000;
	assign font[2][103] = 8'b00000000;
	assign font[3][103] = 8'b00000000;
	assign font[4][103] = 8'b00000000;
	assign font[5][103] = 8'b00000000;
	assign font[6][103] = 8'b00000000;
	assign font[7][103] = 8'b00111100;
	assign font[8][103] = 8'b01000100;
	assign font[9][103] = 8'b01000100;
	assign font[10][103] = 8'b01000100;
	assign font[11][103] = 8'b01000100;
	assign font[12][103] = 8'b01111100;
	assign font[13][103] = 8'b00111100;
	assign font[14][103] = 8'b00000100;
	assign font[15][103] = 8'b00111000;

	assign font[0][104] = 8'b00000000;
	assign font[1][104] = 8'b00000000;
	assign font[2][104] = 8'b00000000;
	assign font[3][104] = 8'b00000000;
	assign font[4][104] = 8'b01100000;
	assign font[5][104] = 8'b01000000;
	assign font[6][104] = 8'b01100000;
	assign font[7][104] = 8'b01011100;
	assign font[8][104] = 8'b01000100;
	assign font[9][104] = 8'b01100100;
	assign font[10][104] = 8'b01100110;
	assign font[11][104] = 8'b01000100;
	assign font[12][104] = 8'b01000100;
	assign font[13][104] = 8'b01100110;
	assign font[14][104] = 8'b00000000;
	assign font[15][104] = 8'b00000000;

	assign font[0][105] = 8'b00000000;
	assign font[1][105] = 8'b00000000;
	assign font[2][105] = 8'b00000000;
	assign font[3][105] = 8'b00000000;
	assign font[4][105] = 8'b00001000;
	assign font[5][105] = 8'b00000000;
	assign font[6][105] = 8'b00000000;
	assign font[7][105] = 8'b00011000;
	assign font[8][105] = 8'b00011000;
	assign font[9][105] = 8'b00001000;
	assign font[10][105] = 8'b00001000;
	assign font[11][105] = 8'b00001000;
	assign font[12][105] = 8'b00001000;
	assign font[13][105] = 8'b00111100;
	assign font[14][105] = 8'b00000000;
	assign font[15][105] = 8'b00000000;

	assign font[0][106] = 8'b00000000;
	assign font[1][106] = 8'b00000000;
	assign font[2][106] = 8'b00000000;
	assign font[3][106] = 8'b00000000;
	assign font[4][106] = 8'b00011000;
	assign font[5][106] = 8'b00000000;
	assign font[6][106] = 8'b00000000;
	assign font[7][106] = 8'b00111000;
	assign font[8][106] = 8'b00011000;
	assign font[9][106] = 8'b00011000;
	assign font[10][106] = 8'b00011000;
	assign font[11][106] = 8'b00011000;
	assign font[12][106] = 8'b00010000;
	assign font[13][106] = 8'b00011000;
	assign font[14][106] = 8'b00010000;
	assign font[15][106] = 8'b01110000;

	assign font[0][107] = 8'b00000000;
	assign font[1][107] = 8'b00000000;
	assign font[2][107] = 8'b00000000;
	assign font[3][107] = 8'b00000000;
	assign font[4][107] = 8'b01000000;
	assign font[5][107] = 8'b01000000;
	assign font[6][107] = 8'b01000000;
	assign font[7][107] = 8'b01001000;
	assign font[8][107] = 8'b01010000;
	assign font[9][107] = 8'b01010000;
	assign font[10][107] = 8'b01110000;
	assign font[11][107] = 8'b01011000;
	assign font[12][107] = 8'b01011000;
	assign font[13][107] = 8'b01001100;
	assign font[14][107] = 8'b00000000;
	assign font[15][107] = 8'b00000000;

	assign font[0][108] = 8'b00000000;
	assign font[1][108] = 8'b00000000;
	assign font[2][108] = 8'b00000000;
	assign font[3][108] = 8'b00000000;
	assign font[4][108] = 8'b00011000;
	assign font[5][108] = 8'b00011000;
	assign font[6][108] = 8'b00011000;
	assign font[7][108] = 8'b00011000;
	assign font[8][108] = 8'b00011000;
	assign font[9][108] = 8'b00011000;
	assign font[10][108] = 8'b00011000;
	assign font[11][108] = 8'b00011000;
	assign font[12][108] = 8'b00011000;
	assign font[13][108] = 8'b00111100;
	assign font[14][108] = 8'b00000000;
	assign font[15][108] = 8'b00000000;

	assign font[0][109] = 8'b00000000;
	assign font[1][109] = 8'b00000000;
	assign font[2][109] = 8'b00000000;
	assign font[3][109] = 8'b00000000;
	assign font[4][109] = 8'b00000000;
	assign font[5][109] = 8'b00000000;
	assign font[6][109] = 8'b00000000;
	assign font[7][109] = 8'b01111100;
	assign font[8][109] = 8'b01110110;
	assign font[9][109] = 8'b01110100;
	assign font[10][109] = 8'b01110110;
	assign font[11][109] = 8'b01110100;
	assign font[12][109] = 8'b01010100;
	assign font[13][109] = 8'b01111110;
	assign font[14][109] = 8'b00000000;
	assign font[15][109] = 8'b00000000;

	assign font[0][110] = 8'b00000000;
	assign font[1][110] = 8'b00000000;
	assign font[2][110] = 8'b00000000;
	assign font[3][110] = 8'b00000000;
	assign font[4][110] = 8'b00000000;
	assign font[5][110] = 8'b00000000;
	assign font[6][110] = 8'b00000000;
	assign font[7][110] = 8'b01111100;
	assign font[8][110] = 8'b01100100;
	assign font[9][110] = 8'b01100110;
	assign font[10][110] = 8'b01000110;
	assign font[11][110] = 8'b01000100;
	assign font[12][110] = 8'b01000100;
	assign font[13][110] = 8'b01100110;
	assign font[14][110] = 8'b00000000;
	assign font[15][110] = 8'b00000000;

	assign font[0][111] = 8'b00000000;
	assign font[1][111] = 8'b00000000;
	assign font[2][111] = 8'b00000000;
	assign font[3][111] = 8'b00000000;
	assign font[4][111] = 8'b00000000;
	assign font[5][111] = 8'b00000000;
	assign font[6][111] = 8'b00000000;
	assign font[7][111] = 8'b00111000;
	assign font[8][111] = 8'b01001000;
	assign font[9][111] = 8'b01001100;
	assign font[10][111] = 8'b01000100;
	assign font[11][111] = 8'b01001100;
	assign font[12][111] = 8'b01001100;
	assign font[13][111] = 8'b00111000;
	assign font[14][111] = 8'b00000000;
	assign font[15][111] = 8'b00000000;

	assign font[0][112] = 8'b00000000;
	assign font[1][112] = 8'b00000000;
	assign font[2][112] = 8'b00000000;
	assign font[3][112] = 8'b00000000;
	assign font[4][112] = 8'b00000000;
	assign font[5][112] = 8'b00000000;
	assign font[6][112] = 8'b00000000;
	assign font[7][112] = 8'b01111000;
	assign font[8][112] = 8'b01101100;
	assign font[9][112] = 8'b01000100;
	assign font[10][112] = 8'b01000100;
	assign font[11][112] = 8'b01001100;
	assign font[12][112] = 8'b01001000;
	assign font[13][112] = 8'b01111000;
	assign font[14][112] = 8'b01000000;
	assign font[15][112] = 8'b01000000;

	assign font[0][113] = 8'b00000000;
	assign font[1][113] = 8'b00000000;
	assign font[2][113] = 8'b00000000;
	assign font[3][113] = 8'b00000000;
	assign font[4][113] = 8'b00000000;
	assign font[5][113] = 8'b00000000;
	assign font[6][113] = 8'b00000000;
	assign font[7][113] = 8'b00111100;
	assign font[8][113] = 8'b01000100;
	assign font[9][113] = 8'b01000100;
	assign font[10][113] = 8'b01000100;
	assign font[11][113] = 8'b01000100;
	assign font[12][113] = 8'b01000100;
	assign font[13][113] = 8'b00111100;
	assign font[14][113] = 8'b00000100;
	assign font[15][113] = 8'b00000100;

	assign font[0][114] = 8'b00000000;
	assign font[1][114] = 8'b00000000;
	assign font[2][114] = 8'b00000000;
	assign font[3][114] = 8'b00000000;
	assign font[4][114] = 8'b00000000;
	assign font[5][114] = 8'b00000000;
	assign font[6][114] = 8'b00000000;
	assign font[7][114] = 8'b01111100;
	assign font[8][114] = 8'b00110110;
	assign font[9][114] = 8'b00100000;
	assign font[10][114] = 8'b00100000;
	assign font[11][114] = 8'b00100000;
	assign font[12][114] = 8'b00100000;
	assign font[13][114] = 8'b01110000;
	assign font[14][114] = 8'b00000000;
	assign font[15][114] = 8'b00000000;

	assign font[0][115] = 8'b00000000;
	assign font[1][115] = 8'b00000000;
	assign font[2][115] = 8'b00000000;
	assign font[3][115] = 8'b00000000;
	assign font[4][115] = 8'b00000000;
	assign font[5][115] = 8'b00000000;
	assign font[6][115] = 8'b00000000;
	assign font[7][115] = 8'b00111000;
	assign font[8][115] = 8'b01000000;
	assign font[9][115] = 8'b01000000;
	assign font[10][115] = 8'b00111000;
	assign font[11][115] = 8'b00111000;
	assign font[12][115] = 8'b00001100;
	assign font[13][115] = 8'b00111000;
	assign font[14][115] = 8'b00000000;
	assign font[15][115] = 8'b00000000;

	assign font[0][116] = 8'b00000000;
	assign font[1][116] = 8'b00000000;
	assign font[2][116] = 8'b00000000;
	assign font[3][116] = 8'b00000000;
	assign font[4][116] = 8'b00110000;
	assign font[5][116] = 8'b00010000;
	assign font[6][116] = 8'b00110000;
	assign font[7][116] = 8'b01111100;
	assign font[8][116] = 8'b00110000;
	assign font[9][116] = 8'b00010000;
	assign font[10][116] = 8'b00010000;
	assign font[11][116] = 8'b00110000;
	assign font[12][116] = 8'b00010000;
	assign font[13][116] = 8'b00011100;
	assign font[14][116] = 8'b00000000;
	assign font[15][116] = 8'b00000000;

	assign font[0][117] = 8'b00000000;
	assign font[1][117] = 8'b00000000;
	assign font[2][117] = 8'b00000000;
	assign font[3][117] = 8'b00000000;
	assign font[4][117] = 8'b00000000;
	assign font[5][117] = 8'b00000000;
	assign font[6][117] = 8'b00000000;
	assign font[7][117] = 8'b01100110;
	assign font[8][117] = 8'b01100100;
	assign font[9][117] = 8'b01100100;
	assign font[10][117] = 8'b01100100;
	assign font[11][117] = 8'b01100100;
	assign font[12][117] = 8'b00100100;
	assign font[13][117] = 8'b00111110;
	assign font[14][117] = 8'b00000000;
	assign font[15][117] = 8'b00000000;

	assign font[0][118] = 8'b00000000;
	assign font[1][118] = 8'b00000000;
	assign font[2][118] = 8'b00000000;
	assign font[3][118] = 8'b00000000;
	assign font[4][118] = 8'b00000000;
	assign font[5][118] = 8'b00000000;
	assign font[6][118] = 8'b00000000;
	assign font[7][118] = 8'b01101100;
	assign font[8][118] = 8'b00101000;
	assign font[9][118] = 8'b00101000;
	assign font[10][118] = 8'b00111000;
	assign font[11][118] = 8'b00010000;
	assign font[12][118] = 8'b00111000;
	assign font[13][118] = 8'b00010000;
	assign font[14][118] = 8'b00000000;
	assign font[15][118] = 8'b00000000;

	assign font[0][119] = 8'b00000000;
	assign font[1][119] = 8'b00000000;
	assign font[2][119] = 8'b00000000;
	assign font[3][119] = 8'b00000000;
	assign font[4][119] = 8'b00000000;
	assign font[5][119] = 8'b00000000;
	assign font[6][119] = 8'b00000000;
	assign font[7][119] = 8'b01111110;
	assign font[8][119] = 8'b01110100;
	assign font[9][119] = 8'b01010100;
	assign font[10][119] = 8'b01011100;
	assign font[11][119] = 8'b01011100;
	assign font[12][119] = 8'b00101000;
	assign font[13][119] = 8'b00101000;
	assign font[14][119] = 8'b00000000;
	assign font[15][119] = 8'b00000000;

	assign font[0][120] = 8'b00000000;
	assign font[1][120] = 8'b00000000;
	assign font[2][120] = 8'b00000000;
	assign font[3][120] = 8'b00000000;
	assign font[4][120] = 8'b00000000;
	assign font[5][120] = 8'b00000000;
	assign font[6][120] = 8'b00000000;
	assign font[7][120] = 8'b00100100;
	assign font[8][120] = 8'b00101100;
	assign font[9][120] = 8'b00101000;
	assign font[10][120] = 8'b00011000;
	assign font[11][120] = 8'b00101000;
	assign font[12][120] = 8'b00101100;
	assign font[13][120] = 8'b00100100;
	assign font[14][120] = 8'b00000000;
	assign font[15][120] = 8'b00000000;

	assign font[0][121] = 8'b00000000;
	assign font[1][121] = 8'b00000000;
	assign font[2][121] = 8'b00000000;
	assign font[3][121] = 8'b00000000;
	assign font[4][121] = 8'b00000000;
	assign font[5][121] = 8'b00000000;
	assign font[6][121] = 8'b00000000;
	assign font[7][121] = 8'b11001100;
	assign font[8][121] = 8'b01101000;
	assign font[9][121] = 8'b01101000;
	assign font[10][121] = 8'b01101000;
	assign font[11][121] = 8'b00111000;
	assign font[12][121] = 8'b00110000;
	assign font[13][121] = 8'b00110000;
	assign font[14][121] = 8'b00100000;
	assign font[15][121] = 8'b01100000;

	assign font[0][122] = 8'b00000000;
	assign font[1][122] = 8'b00000000;
	assign font[2][122] = 8'b00000000;
	assign font[3][122] = 8'b00000000;
	assign font[4][122] = 8'b00000000;
	assign font[5][122] = 8'b00000000;
	assign font[6][122] = 8'b00000000;
	assign font[7][122] = 8'b01111000;
	assign font[8][122] = 8'b00001000;
	assign font[9][122] = 8'b00001000;
	assign font[10][122] = 8'b00010000;
	assign font[11][122] = 8'b01100000;
	assign font[12][122] = 8'b01100000;
	assign font[13][122] = 8'b01111100;
	assign font[14][122] = 8'b00000000;
	assign font[15][122] = 8'b00000000;

	assign font[0][123] = 8'b00000000;
	assign font[1][123] = 8'b00000000;
	assign font[2][123] = 8'b00000000;
	assign font[3][123] = 8'b00000000;
	assign font[4][123] = 8'b00001100;
	assign font[5][123] = 8'b00001000;
	assign font[6][123] = 8'b00010000;
	assign font[7][123] = 8'b00010000;
	assign font[8][123] = 8'b00000000;
	assign font[9][123] = 8'b00100000;
	assign font[10][123] = 8'b00010000;
	assign font[11][123] = 8'b00010000;
	assign font[12][123] = 8'b00010000;
	assign font[13][123] = 8'b00001000;
	assign font[14][123] = 8'b00000100;
	assign font[15][123] = 8'b00000000;

	assign font[0][124] = 8'b00000000;
	assign font[1][124] = 8'b00000000;
	assign font[2][124] = 8'b00000000;
	assign font[3][124] = 8'b00000000;
	assign font[4][124] = 8'b00010000;
	assign font[5][124] = 8'b00010000;
	assign font[6][124] = 8'b00010000;
	assign font[7][124] = 8'b00010000;
	assign font[8][124] = 8'b00010000;
	assign font[9][124] = 8'b00010000;
	assign font[10][124] = 8'b00010000;
	assign font[11][124] = 8'b00010000;
	assign font[12][124] = 8'b00010000;
	assign font[13][124] = 8'b00010000;
	assign font[14][124] = 8'b00010000;
	assign font[15][124] = 8'b00000000;

	assign font[0][125] = 8'b00000000;
	assign font[1][125] = 8'b00000000;
	assign font[2][125] = 8'b00000000;
	assign font[3][125] = 8'b00000000;
	assign font[4][125] = 8'b01100000;
	assign font[5][125] = 8'b00100000;
	assign font[6][125] = 8'b00110000;
	assign font[7][125] = 8'b00110000;
	assign font[8][125] = 8'b00000000;
	assign font[9][125] = 8'b00001000;
	assign font[10][125] = 8'b00110000;
	assign font[11][125] = 8'b00110000;
	assign font[12][125] = 8'b00100000;
	assign font[13][125] = 8'b00100000;
	assign font[14][125] = 8'b01000000;
	assign font[15][125] = 8'b00000000;

	assign font[0][126] = 8'b00000000;
	assign font[1][126] = 8'b00000000;
	assign font[2][126] = 8'b00000000;
	assign font[3][126] = 8'b00000000;
	assign font[4][126] = 8'b00000000;
	assign font[5][126] = 8'b00110110;
	assign font[6][126] = 8'b00110100;
	assign font[7][126] = 8'b00110100;
	assign font[8][126] = 8'b01011100;
	assign font[9][126] = 8'b01001000;
	assign font[10][126] = 8'b00000000;
	assign font[11][126] = 8'b00000000;
	assign font[12][126] = 8'b00000000;
	assign font[13][126] = 8'b00000000;
	assign font[14][126] = 8'b00000000;
	assign font[15][126] = 8'b00000000;

	assign font[0][127] = 8'b11111111;
	assign font[1][127] = 8'b11111111;
	assign font[2][127] = 8'b11111111;
	assign font[3][127] = 8'b11111111;
	assign font[4][127] = 8'b11111111;
	assign font[5][127] = 8'b11111111;
	assign font[6][127] = 8'b11111111;
	assign font[7][127] = 8'b11111111;
	assign font[8][127] = 8'b11111111;
	assign font[9][127] = 8'b11111111;
	assign font[10][127] = 8'b11111111;
	assign font[11][127] = 8'b11111111;
	assign font[12][127] = 8'b11111111;
	assign font[13][127] = 8'b11111111;
	assign font[14][127] = 8'b11111111;
	assign font[15][127] = 8'b11111111;

	assign font[0][128] = 8'b11111111;
	assign font[1][128] = 8'b11111111;
	assign font[2][128] = 8'b11111111;
	assign font[3][128] = 8'b11111111;
	assign font[4][128] = 8'b11111111;
	assign font[5][128] = 8'b11111111;
	assign font[6][128] = 8'b11111111;
	assign font[7][128] = 8'b11111111;
	assign font[8][128] = 8'b11111111;
	assign font[9][128] = 8'b11111111;
	assign font[10][128] = 8'b11111111;
	assign font[11][128] = 8'b11111111;
	assign font[12][128] = 8'b11111111;
	assign font[13][128] = 8'b11111111;
	assign font[14][128] = 8'b11111111;
	assign font[15][128] = 8'b11111111;

	assign font[0][129] = 8'b11111111;
	assign font[1][129] = 8'b11111111;
	assign font[2][129] = 8'b11111111;
	assign font[3][129] = 8'b11111111;
	assign font[4][129] = 8'b11111111;
	assign font[5][129] = 8'b11111111;
	assign font[6][129] = 8'b11111111;
	assign font[7][129] = 8'b11111111;
	assign font[8][129] = 8'b11111111;
	assign font[9][129] = 8'b11111111;
	assign font[10][129] = 8'b11111111;
	assign font[11][129] = 8'b11111111;
	assign font[12][129] = 8'b11111111;
	assign font[13][129] = 8'b11111111;
	assign font[14][129] = 8'b11111111;
	assign font[15][129] = 8'b11111111;

	assign font[0][130] = 8'b11111111;
	assign font[1][130] = 8'b11111111;
	assign font[2][130] = 8'b11111111;
	assign font[3][130] = 8'b11111111;
	assign font[4][130] = 8'b11111111;
	assign font[5][130] = 8'b11111111;
	assign font[6][130] = 8'b11111111;
	assign font[7][130] = 8'b11111111;
	assign font[8][130] = 8'b11111111;
	assign font[9][130] = 8'b11111111;
	assign font[10][130] = 8'b11111111;
	assign font[11][130] = 8'b11111111;
	assign font[12][130] = 8'b11111111;
	assign font[13][130] = 8'b11111111;
	assign font[14][130] = 8'b11111111;
	assign font[15][130] = 8'b11111111;

	assign font[0][131] = 8'b11111111;
	assign font[1][131] = 8'b11111111;
	assign font[2][131] = 8'b11111111;
	assign font[3][131] = 8'b11111111;
	assign font[4][131] = 8'b11111111;
	assign font[5][131] = 8'b11111111;
	assign font[6][131] = 8'b11111111;
	assign font[7][131] = 8'b11111111;
	assign font[8][131] = 8'b11111111;
	assign font[9][131] = 8'b11111111;
	assign font[10][131] = 8'b11111111;
	assign font[11][131] = 8'b11111111;
	assign font[12][131] = 8'b11111111;
	assign font[13][131] = 8'b11111111;
	assign font[14][131] = 8'b11111111;
	assign font[15][131] = 8'b11111111;

	assign font[0][132] = 8'b11111111;
	assign font[1][132] = 8'b11111111;
	assign font[2][132] = 8'b11111111;
	assign font[3][132] = 8'b11111111;
	assign font[4][132] = 8'b11111111;
	assign font[5][132] = 8'b11111111;
	assign font[6][132] = 8'b11111111;
	assign font[7][132] = 8'b11111111;
	assign font[8][132] = 8'b11111111;
	assign font[9][132] = 8'b11111111;
	assign font[10][132] = 8'b11111111;
	assign font[11][132] = 8'b11111111;
	assign font[12][132] = 8'b11111111;
	assign font[13][132] = 8'b11111111;
	assign font[14][132] = 8'b11111111;
	assign font[15][132] = 8'b11111111;

	assign font[0][133] = 8'b11111111;
	assign font[1][133] = 8'b11111111;
	assign font[2][133] = 8'b11111111;
	assign font[3][133] = 8'b11111111;
	assign font[4][133] = 8'b11111111;
	assign font[5][133] = 8'b11111111;
	assign font[6][133] = 8'b11111111;
	assign font[7][133] = 8'b11111111;
	assign font[8][133] = 8'b11111111;
	assign font[9][133] = 8'b11111111;
	assign font[10][133] = 8'b11111111;
	assign font[11][133] = 8'b11111111;
	assign font[12][133] = 8'b11111111;
	assign font[13][133] = 8'b11111111;
	assign font[14][133] = 8'b11111111;
	assign font[15][133] = 8'b11111111;

	assign font[0][134] = 8'b11111111;
	assign font[1][134] = 8'b11111111;
	assign font[2][134] = 8'b11111111;
	assign font[3][134] = 8'b11111111;
	assign font[4][134] = 8'b11111111;
	assign font[5][134] = 8'b11111111;
	assign font[6][134] = 8'b11111111;
	assign font[7][134] = 8'b11111111;
	assign font[8][134] = 8'b11111111;
	assign font[9][134] = 8'b11111111;
	assign font[10][134] = 8'b11111111;
	assign font[11][134] = 8'b11111111;
	assign font[12][134] = 8'b11111111;
	assign font[13][134] = 8'b11111111;
	assign font[14][134] = 8'b11111111;
	assign font[15][134] = 8'b11111111;

	assign font[0][135] = 8'b11111111;
	assign font[1][135] = 8'b11111111;
	assign font[2][135] = 8'b11111111;
	assign font[3][135] = 8'b11111111;
	assign font[4][135] = 8'b11111111;
	assign font[5][135] = 8'b11111111;
	assign font[6][135] = 8'b11111111;
	assign font[7][135] = 8'b11111111;
	assign font[8][135] = 8'b11111111;
	assign font[9][135] = 8'b11111111;
	assign font[10][135] = 8'b11111111;
	assign font[11][135] = 8'b11111111;
	assign font[12][135] = 8'b11111111;
	assign font[13][135] = 8'b11111111;
	assign font[14][135] = 8'b11111111;
	assign font[15][135] = 8'b11111111;

	assign font[0][136] = 8'b11111111;
	assign font[1][136] = 8'b11111111;
	assign font[2][136] = 8'b11111111;
	assign font[3][136] = 8'b11111111;
	assign font[4][136] = 8'b11111111;
	assign font[5][136] = 8'b11111111;
	assign font[6][136] = 8'b11111111;
	assign font[7][136] = 8'b11111111;
	assign font[8][136] = 8'b11111111;
	assign font[9][136] = 8'b11111111;
	assign font[10][136] = 8'b11111111;
	assign font[11][136] = 8'b11111111;
	assign font[12][136] = 8'b11111111;
	assign font[13][136] = 8'b11111111;
	assign font[14][136] = 8'b11111111;
	assign font[15][136] = 8'b11111111;

	assign font[0][137] = 8'b11111111;
	assign font[1][137] = 8'b11111111;
	assign font[2][137] = 8'b11111111;
	assign font[3][137] = 8'b11111111;
	assign font[4][137] = 8'b11111111;
	assign font[5][137] = 8'b11111111;
	assign font[6][137] = 8'b11111111;
	assign font[7][137] = 8'b11111111;
	assign font[8][137] = 8'b11111111;
	assign font[9][137] = 8'b11111111;
	assign font[10][137] = 8'b11111111;
	assign font[11][137] = 8'b11111111;
	assign font[12][137] = 8'b11111111;
	assign font[13][137] = 8'b11111111;
	assign font[14][137] = 8'b11111111;
	assign font[15][137] = 8'b11111111;

	assign font[0][138] = 8'b11111111;
	assign font[1][138] = 8'b11111111;
	assign font[2][138] = 8'b11111111;
	assign font[3][138] = 8'b11111111;
	assign font[4][138] = 8'b11111111;
	assign font[5][138] = 8'b11111111;
	assign font[6][138] = 8'b11111111;
	assign font[7][138] = 8'b11111111;
	assign font[8][138] = 8'b11111111;
	assign font[9][138] = 8'b11111111;
	assign font[10][138] = 8'b11111111;
	assign font[11][138] = 8'b11111111;
	assign font[12][138] = 8'b11111111;
	assign font[13][138] = 8'b11111111;
	assign font[14][138] = 8'b11111111;
	assign font[15][138] = 8'b11111111;

	assign font[0][139] = 8'b11111111;
	assign font[1][139] = 8'b11111111;
	assign font[2][139] = 8'b11111111;
	assign font[3][139] = 8'b11111111;
	assign font[4][139] = 8'b11111111;
	assign font[5][139] = 8'b11111111;
	assign font[6][139] = 8'b11111111;
	assign font[7][139] = 8'b11111111;
	assign font[8][139] = 8'b11111111;
	assign font[9][139] = 8'b11111111;
	assign font[10][139] = 8'b11111111;
	assign font[11][139] = 8'b11111111;
	assign font[12][139] = 8'b11111111;
	assign font[13][139] = 8'b11111111;
	assign font[14][139] = 8'b11111111;
	assign font[15][139] = 8'b11111111;

	assign font[0][140] = 8'b11111111;
	assign font[1][140] = 8'b11111111;
	assign font[2][140] = 8'b11111111;
	assign font[3][140] = 8'b11111111;
	assign font[4][140] = 8'b11111111;
	assign font[5][140] = 8'b11111111;
	assign font[6][140] = 8'b11111111;
	assign font[7][140] = 8'b11111111;
	assign font[8][140] = 8'b11111111;
	assign font[9][140] = 8'b11111111;
	assign font[10][140] = 8'b11111111;
	assign font[11][140] = 8'b11111111;
	assign font[12][140] = 8'b11111111;
	assign font[13][140] = 8'b11111111;
	assign font[14][140] = 8'b11111111;
	assign font[15][140] = 8'b11111111;

	assign font[0][141] = 8'b11111111;
	assign font[1][141] = 8'b11111111;
	assign font[2][141] = 8'b11111111;
	assign font[3][141] = 8'b11111111;
	assign font[4][141] = 8'b11111111;
	assign font[5][141] = 8'b11111111;
	assign font[6][141] = 8'b11111111;
	assign font[7][141] = 8'b11111111;
	assign font[8][141] = 8'b11111111;
	assign font[9][141] = 8'b11111111;
	assign font[10][141] = 8'b11111111;
	assign font[11][141] = 8'b11111111;
	assign font[12][141] = 8'b11111111;
	assign font[13][141] = 8'b11111111;
	assign font[14][141] = 8'b11111111;
	assign font[15][141] = 8'b11111111;

	assign font[0][142] = 8'b11111111;
	assign font[1][142] = 8'b11111111;
	assign font[2][142] = 8'b11111111;
	assign font[3][142] = 8'b11111111;
	assign font[4][142] = 8'b11111111;
	assign font[5][142] = 8'b11111111;
	assign font[6][142] = 8'b11111111;
	assign font[7][142] = 8'b11111111;
	assign font[8][142] = 8'b11111111;
	assign font[9][142] = 8'b11111111;
	assign font[10][142] = 8'b11111111;
	assign font[11][142] = 8'b11111111;
	assign font[12][142] = 8'b11111111;
	assign font[13][142] = 8'b11111111;
	assign font[14][142] = 8'b11111111;
	assign font[15][142] = 8'b11111111;

	assign font[0][143] = 8'b11111111;
	assign font[1][143] = 8'b11111111;
	assign font[2][143] = 8'b11111111;
	assign font[3][143] = 8'b11111111;
	assign font[4][143] = 8'b11111111;
	assign font[5][143] = 8'b11111111;
	assign font[6][143] = 8'b11111111;
	assign font[7][143] = 8'b11111111;
	assign font[8][143] = 8'b11111111;
	assign font[9][143] = 8'b11111111;
	assign font[10][143] = 8'b11111111;
	assign font[11][143] = 8'b11111111;
	assign font[12][143] = 8'b11111111;
	assign font[13][143] = 8'b11111111;
	assign font[14][143] = 8'b11111111;
	assign font[15][143] = 8'b11111111;

	assign font[0][144] = 8'b11111111;
	assign font[1][144] = 8'b11111111;
	assign font[2][144] = 8'b11111111;
	assign font[3][144] = 8'b11111111;
	assign font[4][144] = 8'b11111111;
	assign font[5][144] = 8'b11111111;
	assign font[6][144] = 8'b11111111;
	assign font[7][144] = 8'b11111111;
	assign font[8][144] = 8'b11111111;
	assign font[9][144] = 8'b11111111;
	assign font[10][144] = 8'b11111111;
	assign font[11][144] = 8'b11111111;
	assign font[12][144] = 8'b11111111;
	assign font[13][144] = 8'b11111111;
	assign font[14][144] = 8'b11111111;
	assign font[15][144] = 8'b11111111;

	assign font[0][145] = 8'b11111111;
	assign font[1][145] = 8'b11111111;
	assign font[2][145] = 8'b11111111;
	assign font[3][145] = 8'b11111111;
	assign font[4][145] = 8'b11111111;
	assign font[5][145] = 8'b11111111;
	assign font[6][145] = 8'b11111111;
	assign font[7][145] = 8'b11111111;
	assign font[8][145] = 8'b11111111;
	assign font[9][145] = 8'b11111111;
	assign font[10][145] = 8'b11111111;
	assign font[11][145] = 8'b11111111;
	assign font[12][145] = 8'b11111111;
	assign font[13][145] = 8'b11111111;
	assign font[14][145] = 8'b11111111;
	assign font[15][145] = 8'b11111111;

	assign font[0][146] = 8'b11111111;
	assign font[1][146] = 8'b11111111;
	assign font[2][146] = 8'b11111111;
	assign font[3][146] = 8'b11111111;
	assign font[4][146] = 8'b11111111;
	assign font[5][146] = 8'b11111111;
	assign font[6][146] = 8'b11111111;
	assign font[7][146] = 8'b11111111;
	assign font[8][146] = 8'b11111111;
	assign font[9][146] = 8'b11111111;
	assign font[10][146] = 8'b11111111;
	assign font[11][146] = 8'b11111111;
	assign font[12][146] = 8'b11111111;
	assign font[13][146] = 8'b11111111;
	assign font[14][146] = 8'b11111111;
	assign font[15][146] = 8'b11111111;

	assign font[0][147] = 8'b11111111;
	assign font[1][147] = 8'b11111111;
	assign font[2][147] = 8'b11111111;
	assign font[3][147] = 8'b11111111;
	assign font[4][147] = 8'b11111111;
	assign font[5][147] = 8'b11111111;
	assign font[6][147] = 8'b11111111;
	assign font[7][147] = 8'b11111111;
	assign font[8][147] = 8'b11111111;
	assign font[9][147] = 8'b11111111;
	assign font[10][147] = 8'b11111111;
	assign font[11][147] = 8'b11111111;
	assign font[12][147] = 8'b11111111;
	assign font[13][147] = 8'b11111111;
	assign font[14][147] = 8'b11111111;
	assign font[15][147] = 8'b11111111;

	assign font[0][148] = 8'b11111111;
	assign font[1][148] = 8'b11111111;
	assign font[2][148] = 8'b11111111;
	assign font[3][148] = 8'b11111111;
	assign font[4][148] = 8'b11111111;
	assign font[5][148] = 8'b11111111;
	assign font[6][148] = 8'b11111111;
	assign font[7][148] = 8'b11111111;
	assign font[8][148] = 8'b11111111;
	assign font[9][148] = 8'b11111111;
	assign font[10][148] = 8'b11111111;
	assign font[11][148] = 8'b11111111;
	assign font[12][148] = 8'b11111111;
	assign font[13][148] = 8'b11111111;
	assign font[14][148] = 8'b11111111;
	assign font[15][148] = 8'b11111111;

	assign font[0][149] = 8'b11111111;
	assign font[1][149] = 8'b11111111;
	assign font[2][149] = 8'b11111111;
	assign font[3][149] = 8'b11111111;
	assign font[4][149] = 8'b11111111;
	assign font[5][149] = 8'b11111111;
	assign font[6][149] = 8'b11111111;
	assign font[7][149] = 8'b11111111;
	assign font[8][149] = 8'b11111111;
	assign font[9][149] = 8'b11111111;
	assign font[10][149] = 8'b11111111;
	assign font[11][149] = 8'b11111111;
	assign font[12][149] = 8'b11111111;
	assign font[13][149] = 8'b11111111;
	assign font[14][149] = 8'b11111111;
	assign font[15][149] = 8'b11111111;

	assign font[0][150] = 8'b11111111;
	assign font[1][150] = 8'b11111111;
	assign font[2][150] = 8'b11111111;
	assign font[3][150] = 8'b11111111;
	assign font[4][150] = 8'b11111111;
	assign font[5][150] = 8'b11111111;
	assign font[6][150] = 8'b11111111;
	assign font[7][150] = 8'b11111111;
	assign font[8][150] = 8'b11111111;
	assign font[9][150] = 8'b11111111;
	assign font[10][150] = 8'b11111111;
	assign font[11][150] = 8'b11111111;
	assign font[12][150] = 8'b11111111;
	assign font[13][150] = 8'b11111111;
	assign font[14][150] = 8'b11111111;
	assign font[15][150] = 8'b11111111;

	assign font[0][151] = 8'b11111111;
	assign font[1][151] = 8'b11111111;
	assign font[2][151] = 8'b11111111;
	assign font[3][151] = 8'b11111111;
	assign font[4][151] = 8'b11111111;
	assign font[5][151] = 8'b11111111;
	assign font[6][151] = 8'b11111111;
	assign font[7][151] = 8'b11111111;
	assign font[8][151] = 8'b11111111;
	assign font[9][151] = 8'b11111111;
	assign font[10][151] = 8'b11111111;
	assign font[11][151] = 8'b11111111;
	assign font[12][151] = 8'b11111111;
	assign font[13][151] = 8'b11111111;
	assign font[14][151] = 8'b11111111;
	assign font[15][151] = 8'b11111111;

	assign font[0][152] = 8'b11111111;
	assign font[1][152] = 8'b11111111;
	assign font[2][152] = 8'b11111111;
	assign font[3][152] = 8'b11111111;
	assign font[4][152] = 8'b11111111;
	assign font[5][152] = 8'b11111111;
	assign font[6][152] = 8'b11111111;
	assign font[7][152] = 8'b11111111;
	assign font[8][152] = 8'b11111111;
	assign font[9][152] = 8'b11111111;
	assign font[10][152] = 8'b11111111;
	assign font[11][152] = 8'b11111111;
	assign font[12][152] = 8'b11111111;
	assign font[13][152] = 8'b11111111;
	assign font[14][152] = 8'b11111111;
	assign font[15][152] = 8'b11111111;

	assign font[0][153] = 8'b11111111;
	assign font[1][153] = 8'b11111111;
	assign font[2][153] = 8'b11111111;
	assign font[3][153] = 8'b11111111;
	assign font[4][153] = 8'b11111111;
	assign font[5][153] = 8'b11111111;
	assign font[6][153] = 8'b11111111;
	assign font[7][153] = 8'b11111111;
	assign font[8][153] = 8'b11111111;
	assign font[9][153] = 8'b11111111;
	assign font[10][153] = 8'b11111111;
	assign font[11][153] = 8'b11111111;
	assign font[12][153] = 8'b11111111;
	assign font[13][153] = 8'b11111111;
	assign font[14][153] = 8'b11111111;
	assign font[15][153] = 8'b11111111;

	assign font[0][154] = 8'b11111111;
	assign font[1][154] = 8'b11111111;
	assign font[2][154] = 8'b11111111;
	assign font[3][154] = 8'b11111111;
	assign font[4][154] = 8'b11111111;
	assign font[5][154] = 8'b11111111;
	assign font[6][154] = 8'b11111111;
	assign font[7][154] = 8'b11111111;
	assign font[8][154] = 8'b11111111;
	assign font[9][154] = 8'b11111111;
	assign font[10][154] = 8'b11111111;
	assign font[11][154] = 8'b11111111;
	assign font[12][154] = 8'b11111111;
	assign font[13][154] = 8'b11111111;
	assign font[14][154] = 8'b11111111;
	assign font[15][154] = 8'b11111111;

	assign font[0][155] = 8'b11111111;
	assign font[1][155] = 8'b11111111;
	assign font[2][155] = 8'b11111111;
	assign font[3][155] = 8'b11111111;
	assign font[4][155] = 8'b11111111;
	assign font[5][155] = 8'b11111111;
	assign font[6][155] = 8'b11111111;
	assign font[7][155] = 8'b11111111;
	assign font[8][155] = 8'b11111111;
	assign font[9][155] = 8'b11111111;
	assign font[10][155] = 8'b11111111;
	assign font[11][155] = 8'b11111111;
	assign font[12][155] = 8'b11111111;
	assign font[13][155] = 8'b11111111;
	assign font[14][155] = 8'b11111111;
	assign font[15][155] = 8'b11111111;

	assign font[0][156] = 8'b11111111;
	assign font[1][156] = 8'b11111111;
	assign font[2][156] = 8'b11111111;
	assign font[3][156] = 8'b11111111;
	assign font[4][156] = 8'b11111111;
	assign font[5][156] = 8'b11111111;
	assign font[6][156] = 8'b11111111;
	assign font[7][156] = 8'b11111111;
	assign font[8][156] = 8'b11111111;
	assign font[9][156] = 8'b11111111;
	assign font[10][156] = 8'b11111111;
	assign font[11][156] = 8'b11111111;
	assign font[12][156] = 8'b11111111;
	assign font[13][156] = 8'b11111111;
	assign font[14][156] = 8'b11111111;
	assign font[15][156] = 8'b11111111;

	assign font[0][157] = 8'b11111111;
	assign font[1][157] = 8'b11111111;
	assign font[2][157] = 8'b11111111;
	assign font[3][157] = 8'b11111111;
	assign font[4][157] = 8'b11111111;
	assign font[5][157] = 8'b11111111;
	assign font[6][157] = 8'b11111111;
	assign font[7][157] = 8'b11111111;
	assign font[8][157] = 8'b11111111;
	assign font[9][157] = 8'b11111111;
	assign font[10][157] = 8'b11111111;
	assign font[11][157] = 8'b11111111;
	assign font[12][157] = 8'b11111111;
	assign font[13][157] = 8'b11111111;
	assign font[14][157] = 8'b11111111;
	assign font[15][157] = 8'b11111111;

	assign font[0][158] = 8'b11111111;
	assign font[1][158] = 8'b11111111;
	assign font[2][158] = 8'b11111111;
	assign font[3][158] = 8'b11111111;
	assign font[4][158] = 8'b11111111;
	assign font[5][158] = 8'b11111111;
	assign font[6][158] = 8'b11111111;
	assign font[7][158] = 8'b11111111;
	assign font[8][158] = 8'b11111111;
	assign font[9][158] = 8'b11111111;
	assign font[10][158] = 8'b11111111;
	assign font[11][158] = 8'b11111111;
	assign font[12][158] = 8'b11111111;
	assign font[13][158] = 8'b11111111;
	assign font[14][158] = 8'b11111111;
	assign font[15][158] = 8'b11111111;

	assign font[0][159] = 8'b11111111;
	assign font[1][159] = 8'b11111111;
	assign font[2][159] = 8'b11111111;
	assign font[3][159] = 8'b11111111;
	assign font[4][159] = 8'b11111111;
	assign font[5][159] = 8'b11111111;
	assign font[6][159] = 8'b11111111;
	assign font[7][159] = 8'b11111111;
	assign font[8][159] = 8'b11111111;
	assign font[9][159] = 8'b11111111;
	assign font[10][159] = 8'b11111111;
	assign font[11][159] = 8'b11111111;
	assign font[12][159] = 8'b11111111;
	assign font[13][159] = 8'b11111111;
	assign font[14][159] = 8'b11111111;
	assign font[15][159] = 8'b11111111;

	assign font[0][160] = 8'b11111111;
	assign font[1][160] = 8'b11111111;
	assign font[2][160] = 8'b11111111;
	assign font[3][160] = 8'b11111111;
	assign font[4][160] = 8'b11111111;
	assign font[5][160] = 8'b11111111;
	assign font[6][160] = 8'b11111111;
	assign font[7][160] = 8'b11111111;
	assign font[8][160] = 8'b11111111;
	assign font[9][160] = 8'b11111111;
	assign font[10][160] = 8'b11111111;
	assign font[11][160] = 8'b11111111;
	assign font[12][160] = 8'b11111111;
	assign font[13][160] = 8'b11111111;
	assign font[14][160] = 8'b11111111;
	assign font[15][160] = 8'b11111111;

	assign font[0][161] = 8'b11111111;
	assign font[1][161] = 8'b11111111;
	assign font[2][161] = 8'b11111111;
	assign font[3][161] = 8'b11111111;
	assign font[4][161] = 8'b11111111;
	assign font[5][161] = 8'b11111111;
	assign font[6][161] = 8'b11111111;
	assign font[7][161] = 8'b11111111;
	assign font[8][161] = 8'b11111111;
	assign font[9][161] = 8'b11111111;
	assign font[10][161] = 8'b11111111;
	assign font[11][161] = 8'b11111111;
	assign font[12][161] = 8'b11111111;
	assign font[13][161] = 8'b11111111;
	assign font[14][161] = 8'b11111111;
	assign font[15][161] = 8'b11111111;

	assign font[0][162] = 8'b11111111;
	assign font[1][162] = 8'b11111111;
	assign font[2][162] = 8'b11111111;
	assign font[3][162] = 8'b11111111;
	assign font[4][162] = 8'b11111111;
	assign font[5][162] = 8'b11111111;
	assign font[6][162] = 8'b11111111;
	assign font[7][162] = 8'b11111111;
	assign font[8][162] = 8'b11111111;
	assign font[9][162] = 8'b11111111;
	assign font[10][162] = 8'b11111111;
	assign font[11][162] = 8'b11111111;
	assign font[12][162] = 8'b11111111;
	assign font[13][162] = 8'b11111111;
	assign font[14][162] = 8'b11111111;
	assign font[15][162] = 8'b11111111;

	assign font[0][163] = 8'b11111111;
	assign font[1][163] = 8'b11111111;
	assign font[2][163] = 8'b11111111;
	assign font[3][163] = 8'b11111111;
	assign font[4][163] = 8'b11111111;
	assign font[5][163] = 8'b11111111;
	assign font[6][163] = 8'b11111111;
	assign font[7][163] = 8'b11111111;
	assign font[8][163] = 8'b11111111;
	assign font[9][163] = 8'b11111111;
	assign font[10][163] = 8'b11111111;
	assign font[11][163] = 8'b11111111;
	assign font[12][163] = 8'b11111111;
	assign font[13][163] = 8'b11111111;
	assign font[14][163] = 8'b11111111;
	assign font[15][163] = 8'b11111111;

	assign font[0][164] = 8'b11111111;
	assign font[1][164] = 8'b11111111;
	assign font[2][164] = 8'b11111111;
	assign font[3][164] = 8'b11111111;
	assign font[4][164] = 8'b11111111;
	assign font[5][164] = 8'b11111111;
	assign font[6][164] = 8'b11111111;
	assign font[7][164] = 8'b11111111;
	assign font[8][164] = 8'b11111111;
	assign font[9][164] = 8'b11111111;
	assign font[10][164] = 8'b11111111;
	assign font[11][164] = 8'b11111111;
	assign font[12][164] = 8'b11111111;
	assign font[13][164] = 8'b11111111;
	assign font[14][164] = 8'b11111111;
	assign font[15][164] = 8'b11111111;

	assign font[0][165] = 8'b11111111;
	assign font[1][165] = 8'b11111111;
	assign font[2][165] = 8'b11111111;
	assign font[3][165] = 8'b11111111;
	assign font[4][165] = 8'b11111111;
	assign font[5][165] = 8'b11111111;
	assign font[6][165] = 8'b11111111;
	assign font[7][165] = 8'b11111111;
	assign font[8][165] = 8'b11111111;
	assign font[9][165] = 8'b11111111;
	assign font[10][165] = 8'b11111111;
	assign font[11][165] = 8'b11111111;
	assign font[12][165] = 8'b11111111;
	assign font[13][165] = 8'b11111111;
	assign font[14][165] = 8'b11111111;
	assign font[15][165] = 8'b11111111;

	assign font[0][166] = 8'b11111111;
	assign font[1][166] = 8'b11111111;
	assign font[2][166] = 8'b11111111;
	assign font[3][166] = 8'b11111111;
	assign font[4][166] = 8'b11111111;
	assign font[5][166] = 8'b11111111;
	assign font[6][166] = 8'b11111111;
	assign font[7][166] = 8'b11111111;
	assign font[8][166] = 8'b11111111;
	assign font[9][166] = 8'b11111111;
	assign font[10][166] = 8'b11111111;
	assign font[11][166] = 8'b11111111;
	assign font[12][166] = 8'b11111111;
	assign font[13][166] = 8'b11111111;
	assign font[14][166] = 8'b11111111;
	assign font[15][166] = 8'b11111111;

	assign font[0][167] = 8'b11111111;
	assign font[1][167] = 8'b11111111;
	assign font[2][167] = 8'b11111111;
	assign font[3][167] = 8'b11111111;
	assign font[4][167] = 8'b11111111;
	assign font[5][167] = 8'b11111111;
	assign font[6][167] = 8'b11111111;
	assign font[7][167] = 8'b11111111;
	assign font[8][167] = 8'b11111111;
	assign font[9][167] = 8'b11111111;
	assign font[10][167] = 8'b11111111;
	assign font[11][167] = 8'b11111111;
	assign font[12][167] = 8'b11111111;
	assign font[13][167] = 8'b11111111;
	assign font[14][167] = 8'b11111111;
	assign font[15][167] = 8'b11111111;

	assign font[0][168] = 8'b11111111;
	assign font[1][168] = 8'b11111111;
	assign font[2][168] = 8'b11111111;
	assign font[3][168] = 8'b11111111;
	assign font[4][168] = 8'b11111111;
	assign font[5][168] = 8'b11111111;
	assign font[6][168] = 8'b11111111;
	assign font[7][168] = 8'b11111111;
	assign font[8][168] = 8'b11111111;
	assign font[9][168] = 8'b11111111;
	assign font[10][168] = 8'b11111111;
	assign font[11][168] = 8'b11111111;
	assign font[12][168] = 8'b11111111;
	assign font[13][168] = 8'b11111111;
	assign font[14][168] = 8'b11111111;
	assign font[15][168] = 8'b11111111;

	assign font[0][169] = 8'b11111111;
	assign font[1][169] = 8'b11111111;
	assign font[2][169] = 8'b11111111;
	assign font[3][169] = 8'b11111111;
	assign font[4][169] = 8'b11111111;
	assign font[5][169] = 8'b11111111;
	assign font[6][169] = 8'b11111111;
	assign font[7][169] = 8'b11111111;
	assign font[8][169] = 8'b11111111;
	assign font[9][169] = 8'b11111111;
	assign font[10][169] = 8'b11111111;
	assign font[11][169] = 8'b11111111;
	assign font[12][169] = 8'b11111111;
	assign font[13][169] = 8'b11111111;
	assign font[14][169] = 8'b11111111;
	assign font[15][169] = 8'b11111111;

	assign font[0][170] = 8'b11111111;
	assign font[1][170] = 8'b11111111;
	assign font[2][170] = 8'b11111111;
	assign font[3][170] = 8'b11111111;
	assign font[4][170] = 8'b11111111;
	assign font[5][170] = 8'b11111111;
	assign font[6][170] = 8'b11111111;
	assign font[7][170] = 8'b11111111;
	assign font[8][170] = 8'b11111111;
	assign font[9][170] = 8'b11111111;
	assign font[10][170] = 8'b11111111;
	assign font[11][170] = 8'b11111111;
	assign font[12][170] = 8'b11111111;
	assign font[13][170] = 8'b11111111;
	assign font[14][170] = 8'b11111111;
	assign font[15][170] = 8'b11111111;

	assign font[0][171] = 8'b11111111;
	assign font[1][171] = 8'b11111111;
	assign font[2][171] = 8'b11111111;
	assign font[3][171] = 8'b11111111;
	assign font[4][171] = 8'b11111111;
	assign font[5][171] = 8'b11111111;
	assign font[6][171] = 8'b11111111;
	assign font[7][171] = 8'b11111111;
	assign font[8][171] = 8'b11111111;
	assign font[9][171] = 8'b11111111;
	assign font[10][171] = 8'b11111111;
	assign font[11][171] = 8'b11111111;
	assign font[12][171] = 8'b11111111;
	assign font[13][171] = 8'b11111111;
	assign font[14][171] = 8'b11111111;
	assign font[15][171] = 8'b11111111;

	assign font[0][172] = 8'b11111111;
	assign font[1][172] = 8'b11111111;
	assign font[2][172] = 8'b11111111;
	assign font[3][172] = 8'b11111111;
	assign font[4][172] = 8'b11111111;
	assign font[5][172] = 8'b11111111;
	assign font[6][172] = 8'b11111111;
	assign font[7][172] = 8'b11111111;
	assign font[8][172] = 8'b11111111;
	assign font[9][172] = 8'b11111111;
	assign font[10][172] = 8'b11111111;
	assign font[11][172] = 8'b11111111;
	assign font[12][172] = 8'b11111111;
	assign font[13][172] = 8'b11111111;
	assign font[14][172] = 8'b11111111;
	assign font[15][172] = 8'b11111111;

	assign font[0][173] = 8'b11111111;
	assign font[1][173] = 8'b11111111;
	assign font[2][173] = 8'b11111111;
	assign font[3][173] = 8'b11111111;
	assign font[4][173] = 8'b11111111;
	assign font[5][173] = 8'b11111111;
	assign font[6][173] = 8'b11111111;
	assign font[7][173] = 8'b11111111;
	assign font[8][173] = 8'b11111111;
	assign font[9][173] = 8'b11111111;
	assign font[10][173] = 8'b11111111;
	assign font[11][173] = 8'b11111111;
	assign font[12][173] = 8'b11111111;
	assign font[13][173] = 8'b11111111;
	assign font[14][173] = 8'b11111111;
	assign font[15][173] = 8'b11111111;

	assign font[0][174] = 8'b11111111;
	assign font[1][174] = 8'b11111111;
	assign font[2][174] = 8'b11111111;
	assign font[3][174] = 8'b11111111;
	assign font[4][174] = 8'b11111111;
	assign font[5][174] = 8'b11111111;
	assign font[6][174] = 8'b11111111;
	assign font[7][174] = 8'b11111111;
	assign font[8][174] = 8'b11111111;
	assign font[9][174] = 8'b11111111;
	assign font[10][174] = 8'b11111111;
	assign font[11][174] = 8'b11111111;
	assign font[12][174] = 8'b11111111;
	assign font[13][174] = 8'b11111111;
	assign font[14][174] = 8'b11111111;
	assign font[15][174] = 8'b11111111;

	assign font[0][175] = 8'b11111111;
	assign font[1][175] = 8'b11111111;
	assign font[2][175] = 8'b11111111;
	assign font[3][175] = 8'b11111111;
	assign font[4][175] = 8'b11111111;
	assign font[5][175] = 8'b11111111;
	assign font[6][175] = 8'b11111111;
	assign font[7][175] = 8'b11111111;
	assign font[8][175] = 8'b11111111;
	assign font[9][175] = 8'b11111111;
	assign font[10][175] = 8'b11111111;
	assign font[11][175] = 8'b11111111;
	assign font[12][175] = 8'b11111111;
	assign font[13][175] = 8'b11111111;
	assign font[14][175] = 8'b11111111;
	assign font[15][175] = 8'b11111111;

	assign font[0][176] = 8'b11111111;
	assign font[1][176] = 8'b11111111;
	assign font[2][176] = 8'b11111111;
	assign font[3][176] = 8'b11111111;
	assign font[4][176] = 8'b11111111;
	assign font[5][176] = 8'b11111111;
	assign font[6][176] = 8'b11111111;
	assign font[7][176] = 8'b11111111;
	assign font[8][176] = 8'b11111111;
	assign font[9][176] = 8'b11111111;
	assign font[10][176] = 8'b11111111;
	assign font[11][176] = 8'b11111111;
	assign font[12][176] = 8'b11111111;
	assign font[13][176] = 8'b11111111;
	assign font[14][176] = 8'b11111111;
	assign font[15][176] = 8'b11111111;

	assign font[0][177] = 8'b11111111;
	assign font[1][177] = 8'b11111111;
	assign font[2][177] = 8'b11111111;
	assign font[3][177] = 8'b11111111;
	assign font[4][177] = 8'b11111111;
	assign font[5][177] = 8'b11111111;
	assign font[6][177] = 8'b11111111;
	assign font[7][177] = 8'b11111111;
	assign font[8][177] = 8'b11111111;
	assign font[9][177] = 8'b11111111;
	assign font[10][177] = 8'b11111111;
	assign font[11][177] = 8'b11111111;
	assign font[12][177] = 8'b11111111;
	assign font[13][177] = 8'b11111111;
	assign font[14][177] = 8'b11111111;
	assign font[15][177] = 8'b11111111;

	assign font[0][178] = 8'b11111111;
	assign font[1][178] = 8'b11111111;
	assign font[2][178] = 8'b11111111;
	assign font[3][178] = 8'b11111111;
	assign font[4][178] = 8'b11111111;
	assign font[5][178] = 8'b11111111;
	assign font[6][178] = 8'b11111111;
	assign font[7][178] = 8'b11111111;
	assign font[8][178] = 8'b11111111;
	assign font[9][178] = 8'b11111111;
	assign font[10][178] = 8'b11111111;
	assign font[11][178] = 8'b11111111;
	assign font[12][178] = 8'b11111111;
	assign font[13][178] = 8'b11111111;
	assign font[14][178] = 8'b11111111;
	assign font[15][178] = 8'b11111111;

	assign font[0][179] = 8'b11111111;
	assign font[1][179] = 8'b11111111;
	assign font[2][179] = 8'b11111111;
	assign font[3][179] = 8'b11111111;
	assign font[4][179] = 8'b11111111;
	assign font[5][179] = 8'b11111111;
	assign font[6][179] = 8'b11111111;
	assign font[7][179] = 8'b11111111;
	assign font[8][179] = 8'b11111111;
	assign font[9][179] = 8'b11111111;
	assign font[10][179] = 8'b11111111;
	assign font[11][179] = 8'b11111111;
	assign font[12][179] = 8'b11111111;
	assign font[13][179] = 8'b11111111;
	assign font[14][179] = 8'b11111111;
	assign font[15][179] = 8'b11111111;

	assign font[0][180] = 8'b11111111;
	assign font[1][180] = 8'b11111111;
	assign font[2][180] = 8'b11111111;
	assign font[3][180] = 8'b11111111;
	assign font[4][180] = 8'b11111111;
	assign font[5][180] = 8'b11111111;
	assign font[6][180] = 8'b11111111;
	assign font[7][180] = 8'b11111111;
	assign font[8][180] = 8'b11111111;
	assign font[9][180] = 8'b11111111;
	assign font[10][180] = 8'b11111111;
	assign font[11][180] = 8'b11111111;
	assign font[12][180] = 8'b11111111;
	assign font[13][180] = 8'b11111111;
	assign font[14][180] = 8'b11111111;
	assign font[15][180] = 8'b11111111;

	assign font[0][181] = 8'b11111111;
	assign font[1][181] = 8'b11111111;
	assign font[2][181] = 8'b11111111;
	assign font[3][181] = 8'b11111111;
	assign font[4][181] = 8'b11111111;
	assign font[5][181] = 8'b11111111;
	assign font[6][181] = 8'b11111111;
	assign font[7][181] = 8'b11111111;
	assign font[8][181] = 8'b11111111;
	assign font[9][181] = 8'b11111111;
	assign font[10][181] = 8'b11111111;
	assign font[11][181] = 8'b11111111;
	assign font[12][181] = 8'b11111111;
	assign font[13][181] = 8'b11111111;
	assign font[14][181] = 8'b11111111;
	assign font[15][181] = 8'b11111111;

	assign font[0][182] = 8'b11111111;
	assign font[1][182] = 8'b11111111;
	assign font[2][182] = 8'b11111111;
	assign font[3][182] = 8'b11111111;
	assign font[4][182] = 8'b11111111;
	assign font[5][182] = 8'b11111111;
	assign font[6][182] = 8'b11111111;
	assign font[7][182] = 8'b11111111;
	assign font[8][182] = 8'b11111111;
	assign font[9][182] = 8'b11111111;
	assign font[10][182] = 8'b11111111;
	assign font[11][182] = 8'b11111111;
	assign font[12][182] = 8'b11111111;
	assign font[13][182] = 8'b11111111;
	assign font[14][182] = 8'b11111111;
	assign font[15][182] = 8'b11111111;

	assign font[0][183] = 8'b11111111;
	assign font[1][183] = 8'b11111111;
	assign font[2][183] = 8'b11111111;
	assign font[3][183] = 8'b11111111;
	assign font[4][183] = 8'b11111111;
	assign font[5][183] = 8'b11111111;
	assign font[6][183] = 8'b11111111;
	assign font[7][183] = 8'b11111111;
	assign font[8][183] = 8'b11111111;
	assign font[9][183] = 8'b11111111;
	assign font[10][183] = 8'b11111111;
	assign font[11][183] = 8'b11111111;
	assign font[12][183] = 8'b11111111;
	assign font[13][183] = 8'b11111111;
	assign font[14][183] = 8'b11111111;
	assign font[15][183] = 8'b11111111;

	assign font[0][184] = 8'b11111111;
	assign font[1][184] = 8'b11111111;
	assign font[2][184] = 8'b11111111;
	assign font[3][184] = 8'b11111111;
	assign font[4][184] = 8'b11111111;
	assign font[5][184] = 8'b11111111;
	assign font[6][184] = 8'b11111111;
	assign font[7][184] = 8'b11111111;
	assign font[8][184] = 8'b11111111;
	assign font[9][184] = 8'b11111111;
	assign font[10][184] = 8'b11111111;
	assign font[11][184] = 8'b11111111;
	assign font[12][184] = 8'b11111111;
	assign font[13][184] = 8'b11111111;
	assign font[14][184] = 8'b11111111;
	assign font[15][184] = 8'b11111111;

	assign font[0][185] = 8'b11111111;
	assign font[1][185] = 8'b11111111;
	assign font[2][185] = 8'b11111111;
	assign font[3][185] = 8'b11111111;
	assign font[4][185] = 8'b11111111;
	assign font[5][185] = 8'b11111111;
	assign font[6][185] = 8'b11111111;
	assign font[7][185] = 8'b11111111;
	assign font[8][185] = 8'b11111111;
	assign font[9][185] = 8'b11111111;
	assign font[10][185] = 8'b11111111;
	assign font[11][185] = 8'b11111111;
	assign font[12][185] = 8'b11111111;
	assign font[13][185] = 8'b11111111;
	assign font[14][185] = 8'b11111111;
	assign font[15][185] = 8'b11111111;

	assign font[0][186] = 8'b11111111;
	assign font[1][186] = 8'b11111111;
	assign font[2][186] = 8'b11111111;
	assign font[3][186] = 8'b11111111;
	assign font[4][186] = 8'b11111111;
	assign font[5][186] = 8'b11111111;
	assign font[6][186] = 8'b11111111;
	assign font[7][186] = 8'b11111111;
	assign font[8][186] = 8'b11111111;
	assign font[9][186] = 8'b11111111;
	assign font[10][186] = 8'b11111111;
	assign font[11][186] = 8'b11111111;
	assign font[12][186] = 8'b11111111;
	assign font[13][186] = 8'b11111111;
	assign font[14][186] = 8'b11111111;
	assign font[15][186] = 8'b11111111;

	assign font[0][187] = 8'b11111111;
	assign font[1][187] = 8'b11111111;
	assign font[2][187] = 8'b11111111;
	assign font[3][187] = 8'b11111111;
	assign font[4][187] = 8'b11111111;
	assign font[5][187] = 8'b11111111;
	assign font[6][187] = 8'b11111111;
	assign font[7][187] = 8'b11111111;
	assign font[8][187] = 8'b11111111;
	assign font[9][187] = 8'b11111111;
	assign font[10][187] = 8'b11111111;
	assign font[11][187] = 8'b11111111;
	assign font[12][187] = 8'b11111111;
	assign font[13][187] = 8'b11111111;
	assign font[14][187] = 8'b11111111;
	assign font[15][187] = 8'b11111111;

	assign font[0][188] = 8'b11111111;
	assign font[1][188] = 8'b11111111;
	assign font[2][188] = 8'b11111111;
	assign font[3][188] = 8'b11111111;
	assign font[4][188] = 8'b11111111;
	assign font[5][188] = 8'b11111111;
	assign font[6][188] = 8'b11111111;
	assign font[7][188] = 8'b11111111;
	assign font[8][188] = 8'b11111111;
	assign font[9][188] = 8'b11111111;
	assign font[10][188] = 8'b11111111;
	assign font[11][188] = 8'b11111111;
	assign font[12][188] = 8'b11111111;
	assign font[13][188] = 8'b11111111;
	assign font[14][188] = 8'b11111111;
	assign font[15][188] = 8'b11111111;

	assign font[0][189] = 8'b11111111;
	assign font[1][189] = 8'b11111111;
	assign font[2][189] = 8'b11111111;
	assign font[3][189] = 8'b11111111;
	assign font[4][189] = 8'b11111111;
	assign font[5][189] = 8'b11111111;
	assign font[6][189] = 8'b11111111;
	assign font[7][189] = 8'b11111111;
	assign font[8][189] = 8'b11111111;
	assign font[9][189] = 8'b11111111;
	assign font[10][189] = 8'b11111111;
	assign font[11][189] = 8'b11111111;
	assign font[12][189] = 8'b11111111;
	assign font[13][189] = 8'b11111111;
	assign font[14][189] = 8'b11111111;
	assign font[15][189] = 8'b11111111;

	assign font[0][190] = 8'b11111111;
	assign font[1][190] = 8'b11111111;
	assign font[2][190] = 8'b11111111;
	assign font[3][190] = 8'b11111111;
	assign font[4][190] = 8'b11111111;
	assign font[5][190] = 8'b11111111;
	assign font[6][190] = 8'b11111111;
	assign font[7][190] = 8'b11111111;
	assign font[8][190] = 8'b11111111;
	assign font[9][190] = 8'b11111111;
	assign font[10][190] = 8'b11111111;
	assign font[11][190] = 8'b11111111;
	assign font[12][190] = 8'b11111111;
	assign font[13][190] = 8'b11111111;
	assign font[14][190] = 8'b11111111;
	assign font[15][190] = 8'b11111111;

	assign font[0][191] = 8'b11111111;
	assign font[1][191] = 8'b11111111;
	assign font[2][191] = 8'b11111111;
	assign font[3][191] = 8'b11111111;
	assign font[4][191] = 8'b11111111;
	assign font[5][191] = 8'b11111111;
	assign font[6][191] = 8'b11111111;
	assign font[7][191] = 8'b11111111;
	assign font[8][191] = 8'b11111111;
	assign font[9][191] = 8'b11111111;
	assign font[10][191] = 8'b11111111;
	assign font[11][191] = 8'b11111111;
	assign font[12][191] = 8'b11111111;
	assign font[13][191] = 8'b11111111;
	assign font[14][191] = 8'b11111111;
	assign font[15][191] = 8'b11111111;

	assign font[0][192] = 8'b11111111;
	assign font[1][192] = 8'b11111111;
	assign font[2][192] = 8'b11111111;
	assign font[3][192] = 8'b11111111;
	assign font[4][192] = 8'b11111111;
	assign font[5][192] = 8'b11111111;
	assign font[6][192] = 8'b11111111;
	assign font[7][192] = 8'b11111111;
	assign font[8][192] = 8'b11111111;
	assign font[9][192] = 8'b11111111;
	assign font[10][192] = 8'b11111111;
	assign font[11][192] = 8'b11111111;
	assign font[12][192] = 8'b11111111;
	assign font[13][192] = 8'b11111111;
	assign font[14][192] = 8'b11111111;
	assign font[15][192] = 8'b11111111;

	assign font[0][193] = 8'b11111111;
	assign font[1][193] = 8'b11111111;
	assign font[2][193] = 8'b11111111;
	assign font[3][193] = 8'b11111111;
	assign font[4][193] = 8'b11111111;
	assign font[5][193] = 8'b11111111;
	assign font[6][193] = 8'b11111111;
	assign font[7][193] = 8'b11111111;
	assign font[8][193] = 8'b11111111;
	assign font[9][193] = 8'b11111111;
	assign font[10][193] = 8'b11111111;
	assign font[11][193] = 8'b11111111;
	assign font[12][193] = 8'b11111111;
	assign font[13][193] = 8'b11111111;
	assign font[14][193] = 8'b11111111;
	assign font[15][193] = 8'b11111111;

	assign font[0][194] = 8'b11111111;
	assign font[1][194] = 8'b11111111;
	assign font[2][194] = 8'b11111111;
	assign font[3][194] = 8'b11111111;
	assign font[4][194] = 8'b11111111;
	assign font[5][194] = 8'b11111111;
	assign font[6][194] = 8'b11111111;
	assign font[7][194] = 8'b11111111;
	assign font[8][194] = 8'b11111111;
	assign font[9][194] = 8'b11111111;
	assign font[10][194] = 8'b11111111;
	assign font[11][194] = 8'b11111111;
	assign font[12][194] = 8'b11111111;
	assign font[13][194] = 8'b11111111;
	assign font[14][194] = 8'b11111111;
	assign font[15][194] = 8'b11111111;

	assign font[0][195] = 8'b11111111;
	assign font[1][195] = 8'b11111111;
	assign font[2][195] = 8'b11111111;
	assign font[3][195] = 8'b11111111;
	assign font[4][195] = 8'b11111111;
	assign font[5][195] = 8'b11111111;
	assign font[6][195] = 8'b11111111;
	assign font[7][195] = 8'b11111111;
	assign font[8][195] = 8'b11111111;
	assign font[9][195] = 8'b11111111;
	assign font[10][195] = 8'b11111111;
	assign font[11][195] = 8'b11111111;
	assign font[12][195] = 8'b11111111;
	assign font[13][195] = 8'b11111111;
	assign font[14][195] = 8'b11111111;
	assign font[15][195] = 8'b11111111;

	assign font[0][196] = 8'b11111111;
	assign font[1][196] = 8'b11111111;
	assign font[2][196] = 8'b11111111;
	assign font[3][196] = 8'b11111111;
	assign font[4][196] = 8'b11111111;
	assign font[5][196] = 8'b11111111;
	assign font[6][196] = 8'b11111111;
	assign font[7][196] = 8'b11111111;
	assign font[8][196] = 8'b11111111;
	assign font[9][196] = 8'b11111111;
	assign font[10][196] = 8'b11111111;
	assign font[11][196] = 8'b11111111;
	assign font[12][196] = 8'b11111111;
	assign font[13][196] = 8'b11111111;
	assign font[14][196] = 8'b11111111;
	assign font[15][196] = 8'b11111111;

	assign font[0][197] = 8'b11111111;
	assign font[1][197] = 8'b11111111;
	assign font[2][197] = 8'b11111111;
	assign font[3][197] = 8'b11111111;
	assign font[4][197] = 8'b11111111;
	assign font[5][197] = 8'b11111111;
	assign font[6][197] = 8'b11111111;
	assign font[7][197] = 8'b11111111;
	assign font[8][197] = 8'b11111111;
	assign font[9][197] = 8'b11111111;
	assign font[10][197] = 8'b11111111;
	assign font[11][197] = 8'b11111111;
	assign font[12][197] = 8'b11111111;
	assign font[13][197] = 8'b11111111;
	assign font[14][197] = 8'b11111111;
	assign font[15][197] = 8'b11111111;

	assign font[0][198] = 8'b11111111;
	assign font[1][198] = 8'b11111111;
	assign font[2][198] = 8'b11111111;
	assign font[3][198] = 8'b11111111;
	assign font[4][198] = 8'b11111111;
	assign font[5][198] = 8'b11111111;
	assign font[6][198] = 8'b11111111;
	assign font[7][198] = 8'b11111111;
	assign font[8][198] = 8'b11111111;
	assign font[9][198] = 8'b11111111;
	assign font[10][198] = 8'b11111111;
	assign font[11][198] = 8'b11111111;
	assign font[12][198] = 8'b11111111;
	assign font[13][198] = 8'b11111111;
	assign font[14][198] = 8'b11111111;
	assign font[15][198] = 8'b11111111;

	assign font[0][199] = 8'b11111111;
	assign font[1][199] = 8'b11111111;
	assign font[2][199] = 8'b11111111;
	assign font[3][199] = 8'b11111111;
	assign font[4][199] = 8'b11111111;
	assign font[5][199] = 8'b11111111;
	assign font[6][199] = 8'b11111111;
	assign font[7][199] = 8'b11111111;
	assign font[8][199] = 8'b11111111;
	assign font[9][199] = 8'b11111111;
	assign font[10][199] = 8'b11111111;
	assign font[11][199] = 8'b11111111;
	assign font[12][199] = 8'b11111111;
	assign font[13][199] = 8'b11111111;
	assign font[14][199] = 8'b11111111;
	assign font[15][199] = 8'b11111111;

	assign font[0][200] = 8'b11111111;
	assign font[1][200] = 8'b11111111;
	assign font[2][200] = 8'b11111111;
	assign font[3][200] = 8'b11111111;
	assign font[4][200] = 8'b11111111;
	assign font[5][200] = 8'b11111111;
	assign font[6][200] = 8'b11111111;
	assign font[7][200] = 8'b11111111;
	assign font[8][200] = 8'b11111111;
	assign font[9][200] = 8'b11111111;
	assign font[10][200] = 8'b11111111;
	assign font[11][200] = 8'b11111111;
	assign font[12][200] = 8'b11111111;
	assign font[13][200] = 8'b11111111;
	assign font[14][200] = 8'b11111111;
	assign font[15][200] = 8'b11111111;

	assign font[0][201] = 8'b11111111;
	assign font[1][201] = 8'b11111111;
	assign font[2][201] = 8'b11111111;
	assign font[3][201] = 8'b11111111;
	assign font[4][201] = 8'b11111111;
	assign font[5][201] = 8'b11111111;
	assign font[6][201] = 8'b11111111;
	assign font[7][201] = 8'b11111111;
	assign font[8][201] = 8'b11111111;
	assign font[9][201] = 8'b11111111;
	assign font[10][201] = 8'b11111111;
	assign font[11][201] = 8'b11111111;
	assign font[12][201] = 8'b11111111;
	assign font[13][201] = 8'b11111111;
	assign font[14][201] = 8'b11111111;
	assign font[15][201] = 8'b11111111;

	assign font[0][202] = 8'b11111111;
	assign font[1][202] = 8'b11111111;
	assign font[2][202] = 8'b11111111;
	assign font[3][202] = 8'b11111111;
	assign font[4][202] = 8'b11111111;
	assign font[5][202] = 8'b11111111;
	assign font[6][202] = 8'b11111111;
	assign font[7][202] = 8'b11111111;
	assign font[8][202] = 8'b11111111;
	assign font[9][202] = 8'b11111111;
	assign font[10][202] = 8'b11111111;
	assign font[11][202] = 8'b11111111;
	assign font[12][202] = 8'b11111111;
	assign font[13][202] = 8'b11111111;
	assign font[14][202] = 8'b11111111;
	assign font[15][202] = 8'b11111111;

	assign font[0][203] = 8'b11111111;
	assign font[1][203] = 8'b11111111;
	assign font[2][203] = 8'b11111111;
	assign font[3][203] = 8'b11111111;
	assign font[4][203] = 8'b11111111;
	assign font[5][203] = 8'b11111111;
	assign font[6][203] = 8'b11111111;
	assign font[7][203] = 8'b11111111;
	assign font[8][203] = 8'b11111111;
	assign font[9][203] = 8'b11111111;
	assign font[10][203] = 8'b11111111;
	assign font[11][203] = 8'b11111111;
	assign font[12][203] = 8'b11111111;
	assign font[13][203] = 8'b11111111;
	assign font[14][203] = 8'b11111111;
	assign font[15][203] = 8'b11111111;

	assign font[0][204] = 8'b11111111;
	assign font[1][204] = 8'b11111111;
	assign font[2][204] = 8'b11111111;
	assign font[3][204] = 8'b11111111;
	assign font[4][204] = 8'b11111111;
	assign font[5][204] = 8'b11111111;
	assign font[6][204] = 8'b11111111;
	assign font[7][204] = 8'b11111111;
	assign font[8][204] = 8'b11111111;
	assign font[9][204] = 8'b11111111;
	assign font[10][204] = 8'b11111111;
	assign font[11][204] = 8'b11111111;
	assign font[12][204] = 8'b11111111;
	assign font[13][204] = 8'b11111111;
	assign font[14][204] = 8'b11111111;
	assign font[15][204] = 8'b11111111;

	assign font[0][205] = 8'b11111111;
	assign font[1][205] = 8'b11111111;
	assign font[2][205] = 8'b11111111;
	assign font[3][205] = 8'b11111111;
	assign font[4][205] = 8'b11111111;
	assign font[5][205] = 8'b11111111;
	assign font[6][205] = 8'b11111111;
	assign font[7][205] = 8'b11111111;
	assign font[8][205] = 8'b11111111;
	assign font[9][205] = 8'b11111111;
	assign font[10][205] = 8'b11111111;
	assign font[11][205] = 8'b11111111;
	assign font[12][205] = 8'b11111111;
	assign font[13][205] = 8'b11111111;
	assign font[14][205] = 8'b11111111;
	assign font[15][205] = 8'b11111111;

	assign font[0][206] = 8'b11111111;
	assign font[1][206] = 8'b11111111;
	assign font[2][206] = 8'b11111111;
	assign font[3][206] = 8'b11111111;
	assign font[4][206] = 8'b11111111;
	assign font[5][206] = 8'b11111111;
	assign font[6][206] = 8'b11111111;
	assign font[7][206] = 8'b11111111;
	assign font[8][206] = 8'b11111111;
	assign font[9][206] = 8'b11111111;
	assign font[10][206] = 8'b11111111;
	assign font[11][206] = 8'b11111111;
	assign font[12][206] = 8'b11111111;
	assign font[13][206] = 8'b11111111;
	assign font[14][206] = 8'b11111111;
	assign font[15][206] = 8'b11111111;

	assign font[0][207] = 8'b11111111;
	assign font[1][207] = 8'b11111111;
	assign font[2][207] = 8'b11111111;
	assign font[3][207] = 8'b11111111;
	assign font[4][207] = 8'b11111111;
	assign font[5][207] = 8'b11111111;
	assign font[6][207] = 8'b11111111;
	assign font[7][207] = 8'b11111111;
	assign font[8][207] = 8'b11111111;
	assign font[9][207] = 8'b11111111;
	assign font[10][207] = 8'b11111111;
	assign font[11][207] = 8'b11111111;
	assign font[12][207] = 8'b11111111;
	assign font[13][207] = 8'b11111111;
	assign font[14][207] = 8'b11111111;
	assign font[15][207] = 8'b11111111;

	assign font[0][208] = 8'b11111111;
	assign font[1][208] = 8'b11111111;
	assign font[2][208] = 8'b11111111;
	assign font[3][208] = 8'b11111111;
	assign font[4][208] = 8'b11111111;
	assign font[5][208] = 8'b11111111;
	assign font[6][208] = 8'b11111111;
	assign font[7][208] = 8'b11111111;
	assign font[8][208] = 8'b11111111;
	assign font[9][208] = 8'b11111111;
	assign font[10][208] = 8'b11111111;
	assign font[11][208] = 8'b11111111;
	assign font[12][208] = 8'b11111111;
	assign font[13][208] = 8'b11111111;
	assign font[14][208] = 8'b11111111;
	assign font[15][208] = 8'b11111111;

	assign font[0][209] = 8'b11111111;
	assign font[1][209] = 8'b11111111;
	assign font[2][209] = 8'b11111111;
	assign font[3][209] = 8'b11111111;
	assign font[4][209] = 8'b11111111;
	assign font[5][209] = 8'b11111111;
	assign font[6][209] = 8'b11111111;
	assign font[7][209] = 8'b11111111;
	assign font[8][209] = 8'b11111111;
	assign font[9][209] = 8'b11111111;
	assign font[10][209] = 8'b11111111;
	assign font[11][209] = 8'b11111111;
	assign font[12][209] = 8'b11111111;
	assign font[13][209] = 8'b11111111;
	assign font[14][209] = 8'b11111111;
	assign font[15][209] = 8'b11111111;

	assign font[0][210] = 8'b11111111;
	assign font[1][210] = 8'b11111111;
	assign font[2][210] = 8'b11111111;
	assign font[3][210] = 8'b11111111;
	assign font[4][210] = 8'b11111111;
	assign font[5][210] = 8'b11111111;
	assign font[6][210] = 8'b11111111;
	assign font[7][210] = 8'b11111111;
	assign font[8][210] = 8'b11111111;
	assign font[9][210] = 8'b11111111;
	assign font[10][210] = 8'b11111111;
	assign font[11][210] = 8'b11111111;
	assign font[12][210] = 8'b11111111;
	assign font[13][210] = 8'b11111111;
	assign font[14][210] = 8'b11111111;
	assign font[15][210] = 8'b11111111;

	assign font[0][211] = 8'b11111111;
	assign font[1][211] = 8'b11111111;
	assign font[2][211] = 8'b11111111;
	assign font[3][211] = 8'b11111111;
	assign font[4][211] = 8'b11111111;
	assign font[5][211] = 8'b11111111;
	assign font[6][211] = 8'b11111111;
	assign font[7][211] = 8'b11111111;
	assign font[8][211] = 8'b11111111;
	assign font[9][211] = 8'b11111111;
	assign font[10][211] = 8'b11111111;
	assign font[11][211] = 8'b11111111;
	assign font[12][211] = 8'b11111111;
	assign font[13][211] = 8'b11111111;
	assign font[14][211] = 8'b11111111;
	assign font[15][211] = 8'b11111111;

	assign font[0][212] = 8'b11111111;
	assign font[1][212] = 8'b11111111;
	assign font[2][212] = 8'b11111111;
	assign font[3][212] = 8'b11111111;
	assign font[4][212] = 8'b11111111;
	assign font[5][212] = 8'b11111111;
	assign font[6][212] = 8'b11111111;
	assign font[7][212] = 8'b11111111;
	assign font[8][212] = 8'b11111111;
	assign font[9][212] = 8'b11111111;
	assign font[10][212] = 8'b11111111;
	assign font[11][212] = 8'b11111111;
	assign font[12][212] = 8'b11111111;
	assign font[13][212] = 8'b11111111;
	assign font[14][212] = 8'b11111111;
	assign font[15][212] = 8'b11111111;

	assign font[0][213] = 8'b11111111;
	assign font[1][213] = 8'b11111111;
	assign font[2][213] = 8'b11111111;
	assign font[3][213] = 8'b11111111;
	assign font[4][213] = 8'b11111111;
	assign font[5][213] = 8'b11111111;
	assign font[6][213] = 8'b11111111;
	assign font[7][213] = 8'b11111111;
	assign font[8][213] = 8'b11111111;
	assign font[9][213] = 8'b11111111;
	assign font[10][213] = 8'b11111111;
	assign font[11][213] = 8'b11111111;
	assign font[12][213] = 8'b11111111;
	assign font[13][213] = 8'b11111111;
	assign font[14][213] = 8'b11111111;
	assign font[15][213] = 8'b11111111;

	assign font[0][214] = 8'b11111111;
	assign font[1][214] = 8'b11111111;
	assign font[2][214] = 8'b11111111;
	assign font[3][214] = 8'b11111111;
	assign font[4][214] = 8'b11111111;
	assign font[5][214] = 8'b11111111;
	assign font[6][214] = 8'b11111111;
	assign font[7][214] = 8'b11111111;
	assign font[8][214] = 8'b11111111;
	assign font[9][214] = 8'b11111111;
	assign font[10][214] = 8'b11111111;
	assign font[11][214] = 8'b11111111;
	assign font[12][214] = 8'b11111111;
	assign font[13][214] = 8'b11111111;
	assign font[14][214] = 8'b11111111;
	assign font[15][214] = 8'b11111111;

	assign font[0][215] = 8'b11111111;
	assign font[1][215] = 8'b11111111;
	assign font[2][215] = 8'b11111111;
	assign font[3][215] = 8'b11111111;
	assign font[4][215] = 8'b11111111;
	assign font[5][215] = 8'b11111111;
	assign font[6][215] = 8'b11111111;
	assign font[7][215] = 8'b11111111;
	assign font[8][215] = 8'b11111111;
	assign font[9][215] = 8'b11111111;
	assign font[10][215] = 8'b11111111;
	assign font[11][215] = 8'b11111111;
	assign font[12][215] = 8'b11111111;
	assign font[13][215] = 8'b11111111;
	assign font[14][215] = 8'b11111111;
	assign font[15][215] = 8'b11111111;

	assign font[0][216] = 8'b11111111;
	assign font[1][216] = 8'b11111111;
	assign font[2][216] = 8'b11111111;
	assign font[3][216] = 8'b11111111;
	assign font[4][216] = 8'b11111111;
	assign font[5][216] = 8'b11111111;
	assign font[6][216] = 8'b11111111;
	assign font[7][216] = 8'b11111111;
	assign font[8][216] = 8'b11111111;
	assign font[9][216] = 8'b11111111;
	assign font[10][216] = 8'b11111111;
	assign font[11][216] = 8'b11111111;
	assign font[12][216] = 8'b11111111;
	assign font[13][216] = 8'b11111111;
	assign font[14][216] = 8'b11111111;
	assign font[15][216] = 8'b11111111;

	assign font[0][217] = 8'b11111111;
	assign font[1][217] = 8'b11111111;
	assign font[2][217] = 8'b11111111;
	assign font[3][217] = 8'b11111111;
	assign font[4][217] = 8'b11111111;
	assign font[5][217] = 8'b11111111;
	assign font[6][217] = 8'b11111111;
	assign font[7][217] = 8'b11111111;
	assign font[8][217] = 8'b11111111;
	assign font[9][217] = 8'b11111111;
	assign font[10][217] = 8'b11111111;
	assign font[11][217] = 8'b11111111;
	assign font[12][217] = 8'b11111111;
	assign font[13][217] = 8'b11111111;
	assign font[14][217] = 8'b11111111;
	assign font[15][217] = 8'b11111111;

	assign font[0][218] = 8'b11111111;
	assign font[1][218] = 8'b11111111;
	assign font[2][218] = 8'b11111111;
	assign font[3][218] = 8'b11111111;
	assign font[4][218] = 8'b11111111;
	assign font[5][218] = 8'b11111111;
	assign font[6][218] = 8'b11111111;
	assign font[7][218] = 8'b11111111;
	assign font[8][218] = 8'b11111111;
	assign font[9][218] = 8'b11111111;
	assign font[10][218] = 8'b11111111;
	assign font[11][218] = 8'b11111111;
	assign font[12][218] = 8'b11111111;
	assign font[13][218] = 8'b11111111;
	assign font[14][218] = 8'b11111111;
	assign font[15][218] = 8'b11111111;

	assign font[0][219] = 8'b11111111;
	assign font[1][219] = 8'b11111111;
	assign font[2][219] = 8'b11111111;
	assign font[3][219] = 8'b11111111;
	assign font[4][219] = 8'b11111111;
	assign font[5][219] = 8'b11111111;
	assign font[6][219] = 8'b11111111;
	assign font[7][219] = 8'b11111111;
	assign font[8][219] = 8'b11111111;
	assign font[9][219] = 8'b11111111;
	assign font[10][219] = 8'b11111111;
	assign font[11][219] = 8'b11111111;
	assign font[12][219] = 8'b11111111;
	assign font[13][219] = 8'b11111111;
	assign font[14][219] = 8'b11111111;
	assign font[15][219] = 8'b11111111;

	assign font[0][220] = 8'b11111111;
	assign font[1][220] = 8'b11111111;
	assign font[2][220] = 8'b11111111;
	assign font[3][220] = 8'b11111111;
	assign font[4][220] = 8'b11111111;
	assign font[5][220] = 8'b11111111;
	assign font[6][220] = 8'b11111111;
	assign font[7][220] = 8'b11111111;
	assign font[8][220] = 8'b11111111;
	assign font[9][220] = 8'b11111111;
	assign font[10][220] = 8'b11111111;
	assign font[11][220] = 8'b11111111;
	assign font[12][220] = 8'b11111111;
	assign font[13][220] = 8'b11111111;
	assign font[14][220] = 8'b11111111;
	assign font[15][220] = 8'b11111111;

	assign font[0][221] = 8'b11111111;
	assign font[1][221] = 8'b11111111;
	assign font[2][221] = 8'b11111111;
	assign font[3][221] = 8'b11111111;
	assign font[4][221] = 8'b11111111;
	assign font[5][221] = 8'b11111111;
	assign font[6][221] = 8'b11111111;
	assign font[7][221] = 8'b11111111;
	assign font[8][221] = 8'b11111111;
	assign font[9][221] = 8'b11111111;
	assign font[10][221] = 8'b11111111;
	assign font[11][221] = 8'b11111111;
	assign font[12][221] = 8'b11111111;
	assign font[13][221] = 8'b11111111;
	assign font[14][221] = 8'b11111111;
	assign font[15][221] = 8'b11111111;

	assign font[0][222] = 8'b11111111;
	assign font[1][222] = 8'b11111111;
	assign font[2][222] = 8'b11111111;
	assign font[3][222] = 8'b11111111;
	assign font[4][222] = 8'b11111111;
	assign font[5][222] = 8'b11111111;
	assign font[6][222] = 8'b11111111;
	assign font[7][222] = 8'b11111111;
	assign font[8][222] = 8'b11111111;
	assign font[9][222] = 8'b11111111;
	assign font[10][222] = 8'b11111111;
	assign font[11][222] = 8'b11111111;
	assign font[12][222] = 8'b11111111;
	assign font[13][222] = 8'b11111111;
	assign font[14][222] = 8'b11111111;
	assign font[15][222] = 8'b11111111;

	assign font[0][223] = 8'b11111111;
	assign font[1][223] = 8'b11111111;
	assign font[2][223] = 8'b11111111;
	assign font[3][223] = 8'b11111111;
	assign font[4][223] = 8'b11111111;
	assign font[5][223] = 8'b11111111;
	assign font[6][223] = 8'b11111111;
	assign font[7][223] = 8'b11111111;
	assign font[8][223] = 8'b11111111;
	assign font[9][223] = 8'b11111111;
	assign font[10][223] = 8'b11111111;
	assign font[11][223] = 8'b11111111;
	assign font[12][223] = 8'b11111111;
	assign font[13][223] = 8'b11111111;
	assign font[14][223] = 8'b11111111;
	assign font[15][223] = 8'b11111111;

	assign font[0][224] = 8'b11111111;
	assign font[1][224] = 8'b11111111;
	assign font[2][224] = 8'b11111111;
	assign font[3][224] = 8'b11111111;
	assign font[4][224] = 8'b11111111;
	assign font[5][224] = 8'b11111111;
	assign font[6][224] = 8'b11111111;
	assign font[7][224] = 8'b11111111;
	assign font[8][224] = 8'b11111111;
	assign font[9][224] = 8'b11111111;
	assign font[10][224] = 8'b11111111;
	assign font[11][224] = 8'b11111111;
	assign font[12][224] = 8'b11111111;
	assign font[13][224] = 8'b11111111;
	assign font[14][224] = 8'b11111111;
	assign font[15][224] = 8'b11111111;

	assign font[0][225] = 8'b11111111;
	assign font[1][225] = 8'b11111111;
	assign font[2][225] = 8'b11111111;
	assign font[3][225] = 8'b11111111;
	assign font[4][225] = 8'b11111111;
	assign font[5][225] = 8'b11111111;
	assign font[6][225] = 8'b11111111;
	assign font[7][225] = 8'b11111111;
	assign font[8][225] = 8'b11111111;
	assign font[9][225] = 8'b11111111;
	assign font[10][225] = 8'b11111111;
	assign font[11][225] = 8'b11111111;
	assign font[12][225] = 8'b11111111;
	assign font[13][225] = 8'b11111111;
	assign font[14][225] = 8'b11111111;
	assign font[15][225] = 8'b11111111;

	assign font[0][226] = 8'b11111111;
	assign font[1][226] = 8'b11111111;
	assign font[2][226] = 8'b11111111;
	assign font[3][226] = 8'b11111111;
	assign font[4][226] = 8'b11111111;
	assign font[5][226] = 8'b11111111;
	assign font[6][226] = 8'b11111111;
	assign font[7][226] = 8'b11111111;
	assign font[8][226] = 8'b11111111;
	assign font[9][226] = 8'b11111111;
	assign font[10][226] = 8'b11111111;
	assign font[11][226] = 8'b11111111;
	assign font[12][226] = 8'b11111111;
	assign font[13][226] = 8'b11111111;
	assign font[14][226] = 8'b11111111;
	assign font[15][226] = 8'b11111111;

	assign font[0][227] = 8'b11111111;
	assign font[1][227] = 8'b11111111;
	assign font[2][227] = 8'b11111111;
	assign font[3][227] = 8'b11111111;
	assign font[4][227] = 8'b11111111;
	assign font[5][227] = 8'b11111111;
	assign font[6][227] = 8'b11111111;
	assign font[7][227] = 8'b11111111;
	assign font[8][227] = 8'b11111111;
	assign font[9][227] = 8'b11111111;
	assign font[10][227] = 8'b11111111;
	assign font[11][227] = 8'b11111111;
	assign font[12][227] = 8'b11111111;
	assign font[13][227] = 8'b11111111;
	assign font[14][227] = 8'b11111111;
	assign font[15][227] = 8'b11111111;

	assign font[0][228] = 8'b11111111;
	assign font[1][228] = 8'b11111111;
	assign font[2][228] = 8'b11111111;
	assign font[3][228] = 8'b11111111;
	assign font[4][228] = 8'b11111111;
	assign font[5][228] = 8'b11111111;
	assign font[6][228] = 8'b11111111;
	assign font[7][228] = 8'b11111111;
	assign font[8][228] = 8'b11111111;
	assign font[9][228] = 8'b11111111;
	assign font[10][228] = 8'b11111111;
	assign font[11][228] = 8'b11111111;
	assign font[12][228] = 8'b11111111;
	assign font[13][228] = 8'b11111111;
	assign font[14][228] = 8'b11111111;
	assign font[15][228] = 8'b11111111;

	assign font[0][229] = 8'b11111111;
	assign font[1][229] = 8'b11111111;
	assign font[2][229] = 8'b11111111;
	assign font[3][229] = 8'b11111111;
	assign font[4][229] = 8'b11111111;
	assign font[5][229] = 8'b11111111;
	assign font[6][229] = 8'b11111111;
	assign font[7][229] = 8'b11111111;
	assign font[8][229] = 8'b11111111;
	assign font[9][229] = 8'b11111111;
	assign font[10][229] = 8'b11111111;
	assign font[11][229] = 8'b11111111;
	assign font[12][229] = 8'b11111111;
	assign font[13][229] = 8'b11111111;
	assign font[14][229] = 8'b11111111;
	assign font[15][229] = 8'b11111111;

	assign font[0][230] = 8'b11111111;
	assign font[1][230] = 8'b11111111;
	assign font[2][230] = 8'b11111111;
	assign font[3][230] = 8'b11111111;
	assign font[4][230] = 8'b11111111;
	assign font[5][230] = 8'b11111111;
	assign font[6][230] = 8'b11111111;
	assign font[7][230] = 8'b11111111;
	assign font[8][230] = 8'b11111111;
	assign font[9][230] = 8'b11111111;
	assign font[10][230] = 8'b11111111;
	assign font[11][230] = 8'b11111111;
	assign font[12][230] = 8'b11111111;
	assign font[13][230] = 8'b11111111;
	assign font[14][230] = 8'b11111111;
	assign font[15][230] = 8'b11111111;

	assign font[0][231] = 8'b11111111;
	assign font[1][231] = 8'b11111111;
	assign font[2][231] = 8'b11111111;
	assign font[3][231] = 8'b11111111;
	assign font[4][231] = 8'b11111111;
	assign font[5][231] = 8'b11111111;
	assign font[6][231] = 8'b11111111;
	assign font[7][231] = 8'b11111111;
	assign font[8][231] = 8'b11111111;
	assign font[9][231] = 8'b11111111;
	assign font[10][231] = 8'b11111111;
	assign font[11][231] = 8'b11111111;
	assign font[12][231] = 8'b11111111;
	assign font[13][231] = 8'b11111111;
	assign font[14][231] = 8'b11111111;
	assign font[15][231] = 8'b11111111;

	assign font[0][232] = 8'b11111111;
	assign font[1][232] = 8'b11111111;
	assign font[2][232] = 8'b11111111;
	assign font[3][232] = 8'b11111111;
	assign font[4][232] = 8'b11111111;
	assign font[5][232] = 8'b11111111;
	assign font[6][232] = 8'b11111111;
	assign font[7][232] = 8'b11111111;
	assign font[8][232] = 8'b11111111;
	assign font[9][232] = 8'b11111111;
	assign font[10][232] = 8'b11111111;
	assign font[11][232] = 8'b11111111;
	assign font[12][232] = 8'b11111111;
	assign font[13][232] = 8'b11111111;
	assign font[14][232] = 8'b11111111;
	assign font[15][232] = 8'b11111111;

	assign font[0][233] = 8'b11111111;
	assign font[1][233] = 8'b11111111;
	assign font[2][233] = 8'b11111111;
	assign font[3][233] = 8'b11111111;
	assign font[4][233] = 8'b11111111;
	assign font[5][233] = 8'b11111111;
	assign font[6][233] = 8'b11111111;
	assign font[7][233] = 8'b11111111;
	assign font[8][233] = 8'b11111111;
	assign font[9][233] = 8'b11111111;
	assign font[10][233] = 8'b11111111;
	assign font[11][233] = 8'b11111111;
	assign font[12][233] = 8'b11111111;
	assign font[13][233] = 8'b11111111;
	assign font[14][233] = 8'b11111111;
	assign font[15][233] = 8'b11111111;

	assign font[0][234] = 8'b11111111;
	assign font[1][234] = 8'b11111111;
	assign font[2][234] = 8'b11111111;
	assign font[3][234] = 8'b11111111;
	assign font[4][234] = 8'b11111111;
	assign font[5][234] = 8'b11111111;
	assign font[6][234] = 8'b11111111;
	assign font[7][234] = 8'b11111111;
	assign font[8][234] = 8'b11111111;
	assign font[9][234] = 8'b11111111;
	assign font[10][234] = 8'b11111111;
	assign font[11][234] = 8'b11111111;
	assign font[12][234] = 8'b11111111;
	assign font[13][234] = 8'b11111111;
	assign font[14][234] = 8'b11111111;
	assign font[15][234] = 8'b11111111;

	assign font[0][235] = 8'b11111111;
	assign font[1][235] = 8'b11111111;
	assign font[2][235] = 8'b11111111;
	assign font[3][235] = 8'b11111111;
	assign font[4][235] = 8'b11111111;
	assign font[5][235] = 8'b11111111;
	assign font[6][235] = 8'b11111111;
	assign font[7][235] = 8'b11111111;
	assign font[8][235] = 8'b11111111;
	assign font[9][235] = 8'b11111111;
	assign font[10][235] = 8'b11111111;
	assign font[11][235] = 8'b11111111;
	assign font[12][235] = 8'b11111111;
	assign font[13][235] = 8'b11111111;
	assign font[14][235] = 8'b11111111;
	assign font[15][235] = 8'b11111111;

	assign font[0][236] = 8'b11111111;
	assign font[1][236] = 8'b11111111;
	assign font[2][236] = 8'b11111111;
	assign font[3][236] = 8'b11111111;
	assign font[4][236] = 8'b11111111;
	assign font[5][236] = 8'b11111111;
	assign font[6][236] = 8'b11111111;
	assign font[7][236] = 8'b11111111;
	assign font[8][236] = 8'b11111111;
	assign font[9][236] = 8'b11111111;
	assign font[10][236] = 8'b11111111;
	assign font[11][236] = 8'b11111111;
	assign font[12][236] = 8'b11111111;
	assign font[13][236] = 8'b11111111;
	assign font[14][236] = 8'b11111111;
	assign font[15][236] = 8'b11111111;

	assign font[0][237] = 8'b11111111;
	assign font[1][237] = 8'b11111111;
	assign font[2][237] = 8'b11111111;
	assign font[3][237] = 8'b11111111;
	assign font[4][237] = 8'b11111111;
	assign font[5][237] = 8'b11111111;
	assign font[6][237] = 8'b11111111;
	assign font[7][237] = 8'b11111111;
	assign font[8][237] = 8'b11111111;
	assign font[9][237] = 8'b11111111;
	assign font[10][237] = 8'b11111111;
	assign font[11][237] = 8'b11111111;
	assign font[12][237] = 8'b11111111;
	assign font[13][237] = 8'b11111111;
	assign font[14][237] = 8'b11111111;
	assign font[15][237] = 8'b11111111;

	assign font[0][238] = 8'b11111111;
	assign font[1][238] = 8'b11111111;
	assign font[2][238] = 8'b11111111;
	assign font[3][238] = 8'b11111111;
	assign font[4][238] = 8'b11111111;
	assign font[5][238] = 8'b11111111;
	assign font[6][238] = 8'b11111111;
	assign font[7][238] = 8'b11111111;
	assign font[8][238] = 8'b11111111;
	assign font[9][238] = 8'b11111111;
	assign font[10][238] = 8'b11111111;
	assign font[11][238] = 8'b11111111;
	assign font[12][238] = 8'b11111111;
	assign font[13][238] = 8'b11111111;
	assign font[14][238] = 8'b11111111;
	assign font[15][238] = 8'b11111111;

	assign font[0][239] = 8'b11111111;
	assign font[1][239] = 8'b11111111;
	assign font[2][239] = 8'b11111111;
	assign font[3][239] = 8'b11111111;
	assign font[4][239] = 8'b11111111;
	assign font[5][239] = 8'b11111111;
	assign font[6][239] = 8'b11111111;
	assign font[7][239] = 8'b11111111;
	assign font[8][239] = 8'b11111111;
	assign font[9][239] = 8'b11111111;
	assign font[10][239] = 8'b11111111;
	assign font[11][239] = 8'b11111111;
	assign font[12][239] = 8'b11111111;
	assign font[13][239] = 8'b11111111;
	assign font[14][239] = 8'b11111111;
	assign font[15][239] = 8'b11111111;

	assign font[0][240] = 8'b11111111;
	assign font[1][240] = 8'b11111111;
	assign font[2][240] = 8'b11111111;
	assign font[3][240] = 8'b11111111;
	assign font[4][240] = 8'b11111111;
	assign font[5][240] = 8'b11111111;
	assign font[6][240] = 8'b11111111;
	assign font[7][240] = 8'b11111111;
	assign font[8][240] = 8'b11111111;
	assign font[9][240] = 8'b11111111;
	assign font[10][240] = 8'b11111111;
	assign font[11][240] = 8'b11111111;
	assign font[12][240] = 8'b11111111;
	assign font[13][240] = 8'b11111111;
	assign font[14][240] = 8'b11111111;
	assign font[15][240] = 8'b11111111;

	assign font[0][241] = 8'b11111111;
	assign font[1][241] = 8'b11111111;
	assign font[2][241] = 8'b11111111;
	assign font[3][241] = 8'b11111111;
	assign font[4][241] = 8'b11111111;
	assign font[5][241] = 8'b11111111;
	assign font[6][241] = 8'b11111111;
	assign font[7][241] = 8'b11111111;
	assign font[8][241] = 8'b11111111;
	assign font[9][241] = 8'b11111111;
	assign font[10][241] = 8'b11111111;
	assign font[11][241] = 8'b11111111;
	assign font[12][241] = 8'b11111111;
	assign font[13][241] = 8'b11111111;
	assign font[14][241] = 8'b11111111;
	assign font[15][241] = 8'b11111111;

	assign font[0][242] = 8'b11111111;
	assign font[1][242] = 8'b11111111;
	assign font[2][242] = 8'b11111111;
	assign font[3][242] = 8'b11111111;
	assign font[4][242] = 8'b11111111;
	assign font[5][242] = 8'b11111111;
	assign font[6][242] = 8'b11111111;
	assign font[7][242] = 8'b11111111;
	assign font[8][242] = 8'b11111111;
	assign font[9][242] = 8'b11111111;
	assign font[10][242] = 8'b11111111;
	assign font[11][242] = 8'b11111111;
	assign font[12][242] = 8'b11111111;
	assign font[13][242] = 8'b11111111;
	assign font[14][242] = 8'b11111111;
	assign font[15][242] = 8'b11111111;

	assign font[0][243] = 8'b11111111;
	assign font[1][243] = 8'b11111111;
	assign font[2][243] = 8'b11111111;
	assign font[3][243] = 8'b11111111;
	assign font[4][243] = 8'b11111111;
	assign font[5][243] = 8'b11111111;
	assign font[6][243] = 8'b11111111;
	assign font[7][243] = 8'b11111111;
	assign font[8][243] = 8'b11111111;
	assign font[9][243] = 8'b11111111;
	assign font[10][243] = 8'b11111111;
	assign font[11][243] = 8'b11111111;
	assign font[12][243] = 8'b11111111;
	assign font[13][243] = 8'b11111111;
	assign font[14][243] = 8'b11111111;
	assign font[15][243] = 8'b11111111;

	assign font[0][244] = 8'b11111111;
	assign font[1][244] = 8'b11111111;
	assign font[2][244] = 8'b11111111;
	assign font[3][244] = 8'b11111111;
	assign font[4][244] = 8'b11111111;
	assign font[5][244] = 8'b11111111;
	assign font[6][244] = 8'b11111111;
	assign font[7][244] = 8'b11111111;
	assign font[8][244] = 8'b11111111;
	assign font[9][244] = 8'b11111111;
	assign font[10][244] = 8'b11111111;
	assign font[11][244] = 8'b11111111;
	assign font[12][244] = 8'b11111111;
	assign font[13][244] = 8'b11111111;
	assign font[14][244] = 8'b11111111;
	assign font[15][244] = 8'b11111111;

	assign font[0][245] = 8'b11111111;
	assign font[1][245] = 8'b11111111;
	assign font[2][245] = 8'b11111111;
	assign font[3][245] = 8'b11111111;
	assign font[4][245] = 8'b11111111;
	assign font[5][245] = 8'b11111111;
	assign font[6][245] = 8'b11111111;
	assign font[7][245] = 8'b11111111;
	assign font[8][245] = 8'b11111111;
	assign font[9][245] = 8'b11111111;
	assign font[10][245] = 8'b11111111;
	assign font[11][245] = 8'b11111111;
	assign font[12][245] = 8'b11111111;
	assign font[13][245] = 8'b11111111;
	assign font[14][245] = 8'b11111111;
	assign font[15][245] = 8'b11111111;

	assign font[0][246] = 8'b11111111;
	assign font[1][246] = 8'b11111111;
	assign font[2][246] = 8'b11111111;
	assign font[3][246] = 8'b11111111;
	assign font[4][246] = 8'b11111111;
	assign font[5][246] = 8'b11111111;
	assign font[6][246] = 8'b11111111;
	assign font[7][246] = 8'b11111111;
	assign font[8][246] = 8'b11111111;
	assign font[9][246] = 8'b11111111;
	assign font[10][246] = 8'b11111111;
	assign font[11][246] = 8'b11111111;
	assign font[12][246] = 8'b11111111;
	assign font[13][246] = 8'b11111111;
	assign font[14][246] = 8'b11111111;
	assign font[15][246] = 8'b11111111;

	assign font[0][247] = 8'b11111111;
	assign font[1][247] = 8'b11111111;
	assign font[2][247] = 8'b11111111;
	assign font[3][247] = 8'b11111111;
	assign font[4][247] = 8'b11111111;
	assign font[5][247] = 8'b11111111;
	assign font[6][247] = 8'b11111111;
	assign font[7][247] = 8'b11111111;
	assign font[8][247] = 8'b11111111;
	assign font[9][247] = 8'b11111111;
	assign font[10][247] = 8'b11111111;
	assign font[11][247] = 8'b11111111;
	assign font[12][247] = 8'b11111111;
	assign font[13][247] = 8'b11111111;
	assign font[14][247] = 8'b11111111;
	assign font[15][247] = 8'b11111111;

	assign font[0][248] = 8'b11111111;
	assign font[1][248] = 8'b11111111;
	assign font[2][248] = 8'b11111111;
	assign font[3][248] = 8'b11111111;
	assign font[4][248] = 8'b11111111;
	assign font[5][248] = 8'b11111111;
	assign font[6][248] = 8'b11111111;
	assign font[7][248] = 8'b11111111;
	assign font[8][248] = 8'b11111111;
	assign font[9][248] = 8'b11111111;
	assign font[10][248] = 8'b11111111;
	assign font[11][248] = 8'b11111111;
	assign font[12][248] = 8'b11111111;
	assign font[13][248] = 8'b11111111;
	assign font[14][248] = 8'b11111111;
	assign font[15][248] = 8'b11111111;

	assign font[0][249] = 8'b11111111;
	assign font[1][249] = 8'b11111111;
	assign font[2][249] = 8'b11111111;
	assign font[3][249] = 8'b11111111;
	assign font[4][249] = 8'b11111111;
	assign font[5][249] = 8'b11111111;
	assign font[6][249] = 8'b11111111;
	assign font[7][249] = 8'b11111111;
	assign font[8][249] = 8'b11111111;
	assign font[9][249] = 8'b11111111;
	assign font[10][249] = 8'b11111111;
	assign font[11][249] = 8'b11111111;
	assign font[12][249] = 8'b11111111;
	assign font[13][249] = 8'b11111111;
	assign font[14][249] = 8'b11111111;
	assign font[15][249] = 8'b11111111;

	assign font[0][250] = 8'b11111111;
	assign font[1][250] = 8'b11111111;
	assign font[2][250] = 8'b11111111;
	assign font[3][250] = 8'b11111111;
	assign font[4][250] = 8'b11111111;
	assign font[5][250] = 8'b11111111;
	assign font[6][250] = 8'b11111111;
	assign font[7][250] = 8'b11111111;
	assign font[8][250] = 8'b11111111;
	assign font[9][250] = 8'b11111111;
	assign font[10][250] = 8'b11111111;
	assign font[11][250] = 8'b11111111;
	assign font[12][250] = 8'b11111111;
	assign font[13][250] = 8'b11111111;
	assign font[14][250] = 8'b11111111;
	assign font[15][250] = 8'b11111111;

	assign font[0][251] = 8'b11111111;
	assign font[1][251] = 8'b11111111;
	assign font[2][251] = 8'b11111111;
	assign font[3][251] = 8'b11111111;
	assign font[4][251] = 8'b11111111;
	assign font[5][251] = 8'b11111111;
	assign font[6][251] = 8'b11111111;
	assign font[7][251] = 8'b11111111;
	assign font[8][251] = 8'b11111111;
	assign font[9][251] = 8'b11111111;
	assign font[10][251] = 8'b11111111;
	assign font[11][251] = 8'b11111111;
	assign font[12][251] = 8'b11111111;
	assign font[13][251] = 8'b11111111;
	assign font[14][251] = 8'b11111111;
	assign font[15][251] = 8'b11111111;

	assign font[0][252] = 8'b11111111;
	assign font[1][252] = 8'b11111111;
	assign font[2][252] = 8'b11111111;
	assign font[3][252] = 8'b11111111;
	assign font[4][252] = 8'b11111111;
	assign font[5][252] = 8'b11111111;
	assign font[6][252] = 8'b11111111;
	assign font[7][252] = 8'b11111111;
	assign font[8][252] = 8'b11111111;
	assign font[9][252] = 8'b11111111;
	assign font[10][252] = 8'b11111111;
	assign font[11][252] = 8'b11111111;
	assign font[12][252] = 8'b11111111;
	assign font[13][252] = 8'b11111111;
	assign font[14][252] = 8'b11111111;
	assign font[15][252] = 8'b11111111;

	assign font[0][253] = 8'b11111111;
	assign font[1][253] = 8'b11111111;
	assign font[2][253] = 8'b11111111;
	assign font[3][253] = 8'b11111111;
	assign font[4][253] = 8'b11111111;
	assign font[5][253] = 8'b11111111;
	assign font[6][253] = 8'b11111111;
	assign font[7][253] = 8'b11111111;
	assign font[8][253] = 8'b11111111;
	assign font[9][253] = 8'b11111111;
	assign font[10][253] = 8'b11111111;
	assign font[11][253] = 8'b11111111;
	assign font[12][253] = 8'b11111111;
	assign font[13][253] = 8'b11111111;
	assign font[14][253] = 8'b11111111;
	assign font[15][253] = 8'b11111111;

	assign font[0][254] = 8'b11111111;
	assign font[1][254] = 8'b11111111;
	assign font[2][254] = 8'b11111111;
	assign font[3][254] = 8'b11111111;
	assign font[4][254] = 8'b11111111;
	assign font[5][254] = 8'b11111111;
	assign font[6][254] = 8'b11111111;
	assign font[7][254] = 8'b11111111;
	assign font[8][254] = 8'b11111111;
	assign font[9][254] = 8'b11111111;
	assign font[10][254] = 8'b11111111;
	assign font[11][254] = 8'b11111111;
	assign font[12][254] = 8'b11111111;
	assign font[13][254] = 8'b11111111;
	assign font[14][254] = 8'b11111111;
	assign font[15][254] = 8'b11111111;

	assign font[0][255] = 8'b11111111;
	assign font[1][255] = 8'b11111111;
	assign font[2][255] = 8'b11111111;
	assign font[3][255] = 8'b11111111;
	assign font[4][255] = 8'b11111111;
	assign font[5][255] = 8'b11111111;
	assign font[6][255] = 8'b11111111;
	assign font[7][255] = 8'b11111111;
	assign font[8][255] = 8'b11111111;
	assign font[9][255] = 8'b11111111;
	assign font[10][255] = 8'b11111111;
	assign font[11][255] = 8'b11111111;
	assign font[12][255] = 8'b11111111;
	assign font[13][255] = 8'b11111111;
	assign font[14][255] = 8'b11111111;
	assign font[15][255] = 8'b11111111;



  assign pixel = font[sym_y][sym_code][sym_x];
endmodule

`define FONT_HEIGHT 32
`define FONT_WIDTH  14

module font_vt323_14x32
(
  input wire  [$clog2(`FONT_WIDTH)-1:0]  sym_x,
  input wire  [$clog2(`FONT_HEIGHT)-1:0] sym_y,
  input wire  [7:0]              sym_code,
  output wire                    sym_pixel
);

  wire [0:`FONT_WIDTH-1] font [`FONT_HEIGHT-1:0] [255:0];

// Here all font bits should be assigned
	assign font[0][0] = 14'b11111111111111;
	assign font[1][0] = 14'b11111111111111;
	assign font[2][0] = 14'b11111111111111;
	assign font[3][0] = 14'b11111111111111;
	assign font[4][0] = 14'b11111111111111;
	assign font[5][0] = 14'b11111111111111;
	assign font[6][0] = 14'b11111111111111;
	assign font[7][0] = 14'b11111111111111;
	assign font[8][0] = 14'b11111111111111;
	assign font[9][0] = 14'b11111111111111;
	assign font[10][0] = 14'b11111111111111;
	assign font[11][0] = 14'b11111111111111;
	assign font[12][0] = 14'b11111111111111;
	assign font[13][0] = 14'b11111111111111;
	assign font[14][0] = 14'b11111111111111;
	assign font[15][0] = 14'b11111111111111;
	assign font[16][0] = 14'b11111111111111;
	assign font[17][0] = 14'b11111111111111;
	assign font[18][0] = 14'b11111111111111;
	assign font[19][0] = 14'b11111111111111;
	assign font[20][0] = 14'b11111111111111;
	assign font[21][0] = 14'b11111111111111;
	assign font[22][0] = 14'b11111111111111;
	assign font[23][0] = 14'b11111111111111;
	assign font[24][0] = 14'b11111111111111;
	assign font[25][0] = 14'b11111111111111;
	assign font[26][0] = 14'b11111111111111;
	assign font[27][0] = 14'b11111111111111;
	assign font[28][0] = 14'b11111111111111;
	assign font[29][0] = 14'b11111111111111;
	assign font[30][0] = 14'b11111111111111;
	assign font[31][0] = 14'b11111111111111;

	assign font[0][1] = 14'b11111111111111;
	assign font[1][1] = 14'b11111111111111;
	assign font[2][1] = 14'b11111111111111;
	assign font[3][1] = 14'b11111111111111;
	assign font[4][1] = 14'b11111111111111;
	assign font[5][1] = 14'b11111111111111;
	assign font[6][1] = 14'b11111111111111;
	assign font[7][1] = 14'b11111111111111;
	assign font[8][1] = 14'b11111111111111;
	assign font[9][1] = 14'b11111111111111;
	assign font[10][1] = 14'b11111111111111;
	assign font[11][1] = 14'b11111111111111;
	assign font[12][1] = 14'b11111111111111;
	assign font[13][1] = 14'b11111111111111;
	assign font[14][1] = 14'b11111111111111;
	assign font[15][1] = 14'b11111111111111;
	assign font[16][1] = 14'b11111111111111;
	assign font[17][1] = 14'b11111111111111;
	assign font[18][1] = 14'b11111111111111;
	assign font[19][1] = 14'b11111111111111;
	assign font[20][1] = 14'b11111111111111;
	assign font[21][1] = 14'b11111111111111;
	assign font[22][1] = 14'b11111111111111;
	assign font[23][1] = 14'b11111111111111;
	assign font[24][1] = 14'b11111111111111;
	assign font[25][1] = 14'b11111111111111;
	assign font[26][1] = 14'b11111111111111;
	assign font[27][1] = 14'b11111111111111;
	assign font[28][1] = 14'b11111111111111;
	assign font[29][1] = 14'b11111111111111;
	assign font[30][1] = 14'b11111111111111;
	assign font[31][1] = 14'b11111111111111;

	assign font[0][2] = 14'b11111111111111;
	assign font[1][2] = 14'b11111111111111;
	assign font[2][2] = 14'b11111111111111;
	assign font[3][2] = 14'b11111111111111;
	assign font[4][2] = 14'b11111111111111;
	assign font[5][2] = 14'b11111111111111;
	assign font[6][2] = 14'b11111111111111;
	assign font[7][2] = 14'b11111111111111;
	assign font[8][2] = 14'b11111111111111;
	assign font[9][2] = 14'b11111111111111;
	assign font[10][2] = 14'b11111111111111;
	assign font[11][2] = 14'b11111111111111;
	assign font[12][2] = 14'b11111111111111;
	assign font[13][2] = 14'b11111111111111;
	assign font[14][2] = 14'b11111111111111;
	assign font[15][2] = 14'b11111111111111;
	assign font[16][2] = 14'b11111111111111;
	assign font[17][2] = 14'b11111111111111;
	assign font[18][2] = 14'b11111111111111;
	assign font[19][2] = 14'b11111111111111;
	assign font[20][2] = 14'b11111111111111;
	assign font[21][2] = 14'b11111111111111;
	assign font[22][2] = 14'b11111111111111;
	assign font[23][2] = 14'b11111111111111;
	assign font[24][2] = 14'b11111111111111;
	assign font[25][2] = 14'b11111111111111;
	assign font[26][2] = 14'b11111111111111;
	assign font[27][2] = 14'b11111111111111;
	assign font[28][2] = 14'b11111111111111;
	assign font[29][2] = 14'b11111111111111;
	assign font[30][2] = 14'b11111111111111;
	assign font[31][2] = 14'b11111111111111;

	assign font[0][3] = 14'b11111111111111;
	assign font[1][3] = 14'b11111111111111;
	assign font[2][3] = 14'b11111111111111;
	assign font[3][3] = 14'b11111111111111;
	assign font[4][3] = 14'b11111111111111;
	assign font[5][3] = 14'b11111111111111;
	assign font[6][3] = 14'b11111111111111;
	assign font[7][3] = 14'b11111111111111;
	assign font[8][3] = 14'b11111111111111;
	assign font[9][3] = 14'b11111111111111;
	assign font[10][3] = 14'b11111111111111;
	assign font[11][3] = 14'b11111111111111;
	assign font[12][3] = 14'b11111111111111;
	assign font[13][3] = 14'b11111111111111;
	assign font[14][3] = 14'b11111111111111;
	assign font[15][3] = 14'b11111111111111;
	assign font[16][3] = 14'b11111111111111;
	assign font[17][3] = 14'b11111111111111;
	assign font[18][3] = 14'b11111111111111;
	assign font[19][3] = 14'b11111111111111;
	assign font[20][3] = 14'b11111111111111;
	assign font[21][3] = 14'b11111111111111;
	assign font[22][3] = 14'b11111111111111;
	assign font[23][3] = 14'b11111111111111;
	assign font[24][3] = 14'b11111111111111;
	assign font[25][3] = 14'b11111111111111;
	assign font[26][3] = 14'b11111111111111;
	assign font[27][3] = 14'b11111111111111;
	assign font[28][3] = 14'b11111111111111;
	assign font[29][3] = 14'b11111111111111;
	assign font[30][3] = 14'b11111111111111;
	assign font[31][3] = 14'b11111111111111;

	assign font[0][4] = 14'b11111111111111;
	assign font[1][4] = 14'b11111111111111;
	assign font[2][4] = 14'b11111111111111;
	assign font[3][4] = 14'b11111111111111;
	assign font[4][4] = 14'b11111111111111;
	assign font[5][4] = 14'b11111111111111;
	assign font[6][4] = 14'b11111111111111;
	assign font[7][4] = 14'b11111111111111;
	assign font[8][4] = 14'b11111111111111;
	assign font[9][4] = 14'b11111111111111;
	assign font[10][4] = 14'b11111111111111;
	assign font[11][4] = 14'b11111111111111;
	assign font[12][4] = 14'b11111111111111;
	assign font[13][4] = 14'b11111111111111;
	assign font[14][4] = 14'b11111111111111;
	assign font[15][4] = 14'b11111111111111;
	assign font[16][4] = 14'b11111111111111;
	assign font[17][4] = 14'b11111111111111;
	assign font[18][4] = 14'b11111111111111;
	assign font[19][4] = 14'b11111111111111;
	assign font[20][4] = 14'b11111111111111;
	assign font[21][4] = 14'b11111111111111;
	assign font[22][4] = 14'b11111111111111;
	assign font[23][4] = 14'b11111111111111;
	assign font[24][4] = 14'b11111111111111;
	assign font[25][4] = 14'b11111111111111;
	assign font[26][4] = 14'b11111111111111;
	assign font[27][4] = 14'b11111111111111;
	assign font[28][4] = 14'b11111111111111;
	assign font[29][4] = 14'b11111111111111;
	assign font[30][4] = 14'b11111111111111;
	assign font[31][4] = 14'b11111111111111;

	assign font[0][5] = 14'b11111111111111;
	assign font[1][5] = 14'b11111111111111;
	assign font[2][5] = 14'b11111111111111;
	assign font[3][5] = 14'b11111111111111;
	assign font[4][5] = 14'b11111111111111;
	assign font[5][5] = 14'b11111111111111;
	assign font[6][5] = 14'b11111111111111;
	assign font[7][5] = 14'b11111111111111;
	assign font[8][5] = 14'b11111111111111;
	assign font[9][5] = 14'b11111111111111;
	assign font[10][5] = 14'b11111111111111;
	assign font[11][5] = 14'b11111111111111;
	assign font[12][5] = 14'b11111111111111;
	assign font[13][5] = 14'b11111111111111;
	assign font[14][5] = 14'b11111111111111;
	assign font[15][5] = 14'b11111111111111;
	assign font[16][5] = 14'b11111111111111;
	assign font[17][5] = 14'b11111111111111;
	assign font[18][5] = 14'b11111111111111;
	assign font[19][5] = 14'b11111111111111;
	assign font[20][5] = 14'b11111111111111;
	assign font[21][5] = 14'b11111111111111;
	assign font[22][5] = 14'b11111111111111;
	assign font[23][5] = 14'b11111111111111;
	assign font[24][5] = 14'b11111111111111;
	assign font[25][5] = 14'b11111111111111;
	assign font[26][5] = 14'b11111111111111;
	assign font[27][5] = 14'b11111111111111;
	assign font[28][5] = 14'b11111111111111;
	assign font[29][5] = 14'b11111111111111;
	assign font[30][5] = 14'b11111111111111;
	assign font[31][5] = 14'b11111111111111;

	assign font[0][6] = 14'b11111111111111;
	assign font[1][6] = 14'b11111111111111;
	assign font[2][6] = 14'b11111111111111;
	assign font[3][6] = 14'b11111111111111;
	assign font[4][6] = 14'b11111111111111;
	assign font[5][6] = 14'b11111111111111;
	assign font[6][6] = 14'b11111111111111;
	assign font[7][6] = 14'b11111111111111;
	assign font[8][6] = 14'b11111111111111;
	assign font[9][6] = 14'b11111111111111;
	assign font[10][6] = 14'b11111111111111;
	assign font[11][6] = 14'b11111111111111;
	assign font[12][6] = 14'b11111111111111;
	assign font[13][6] = 14'b11111111111111;
	assign font[14][6] = 14'b11111111111111;
	assign font[15][6] = 14'b11111111111111;
	assign font[16][6] = 14'b11111111111111;
	assign font[17][6] = 14'b11111111111111;
	assign font[18][6] = 14'b11111111111111;
	assign font[19][6] = 14'b11111111111111;
	assign font[20][6] = 14'b11111111111111;
	assign font[21][6] = 14'b11111111111111;
	assign font[22][6] = 14'b11111111111111;
	assign font[23][6] = 14'b11111111111111;
	assign font[24][6] = 14'b11111111111111;
	assign font[25][6] = 14'b11111111111111;
	assign font[26][6] = 14'b11111111111111;
	assign font[27][6] = 14'b11111111111111;
	assign font[28][6] = 14'b11111111111111;
	assign font[29][6] = 14'b11111111111111;
	assign font[30][6] = 14'b11111111111111;
	assign font[31][6] = 14'b11111111111111;

	assign font[0][7] = 14'b11111111111111;
	assign font[1][7] = 14'b11111111111111;
	assign font[2][7] = 14'b11111111111111;
	assign font[3][7] = 14'b11111111111111;
	assign font[4][7] = 14'b11111111111111;
	assign font[5][7] = 14'b11111111111111;
	assign font[6][7] = 14'b11111111111111;
	assign font[7][7] = 14'b11111111111111;
	assign font[8][7] = 14'b11111111111111;
	assign font[9][7] = 14'b11111111111111;
	assign font[10][7] = 14'b11111111111111;
	assign font[11][7] = 14'b11111111111111;
	assign font[12][7] = 14'b11111111111111;
	assign font[13][7] = 14'b11111111111111;
	assign font[14][7] = 14'b11111111111111;
	assign font[15][7] = 14'b11111111111111;
	assign font[16][7] = 14'b11111111111111;
	assign font[17][7] = 14'b11111111111111;
	assign font[18][7] = 14'b11111111111111;
	assign font[19][7] = 14'b11111111111111;
	assign font[20][7] = 14'b11111111111111;
	assign font[21][7] = 14'b11111111111111;
	assign font[22][7] = 14'b11111111111111;
	assign font[23][7] = 14'b11111111111111;
	assign font[24][7] = 14'b11111111111111;
	assign font[25][7] = 14'b11111111111111;
	assign font[26][7] = 14'b11111111111111;
	assign font[27][7] = 14'b11111111111111;
	assign font[28][7] = 14'b11111111111111;
	assign font[29][7] = 14'b11111111111111;
	assign font[30][7] = 14'b11111111111111;
	assign font[31][7] = 14'b11111111111111;

	assign font[0][8] = 14'b11111111111111;
	assign font[1][8] = 14'b11111111111111;
	assign font[2][8] = 14'b11111111111111;
	assign font[3][8] = 14'b11111111111111;
	assign font[4][8] = 14'b11111111111111;
	assign font[5][8] = 14'b11111111111111;
	assign font[6][8] = 14'b11111111111111;
	assign font[7][8] = 14'b11111111111111;
	assign font[8][8] = 14'b11111111111111;
	assign font[9][8] = 14'b11111111111111;
	assign font[10][8] = 14'b11111111111111;
	assign font[11][8] = 14'b11111111111111;
	assign font[12][8] = 14'b11111111111111;
	assign font[13][8] = 14'b11111111111111;
	assign font[14][8] = 14'b11111111111111;
	assign font[15][8] = 14'b11111111111111;
	assign font[16][8] = 14'b11111111111111;
	assign font[17][8] = 14'b11111111111111;
	assign font[18][8] = 14'b11111111111111;
	assign font[19][8] = 14'b11111111111111;
	assign font[20][8] = 14'b11111111111111;
	assign font[21][8] = 14'b11111111111111;
	assign font[22][8] = 14'b11111111111111;
	assign font[23][8] = 14'b11111111111111;
	assign font[24][8] = 14'b11111111111111;
	assign font[25][8] = 14'b11111111111111;
	assign font[26][8] = 14'b11111111111111;
	assign font[27][8] = 14'b11111111111111;
	assign font[28][8] = 14'b11111111111111;
	assign font[29][8] = 14'b11111111111111;
	assign font[30][8] = 14'b11111111111111;
	assign font[31][8] = 14'b11111111111111;

	assign font[0][9] = 14'b11111111111111;
	assign font[1][9] = 14'b11111111111111;
	assign font[2][9] = 14'b11111111111111;
	assign font[3][9] = 14'b11111111111111;
	assign font[4][9] = 14'b11111111111111;
	assign font[5][9] = 14'b11111111111111;
	assign font[6][9] = 14'b11111111111111;
	assign font[7][9] = 14'b11111111111111;
	assign font[8][9] = 14'b11111111111111;
	assign font[9][9] = 14'b11111111111111;
	assign font[10][9] = 14'b11111111111111;
	assign font[11][9] = 14'b11111111111111;
	assign font[12][9] = 14'b11111111111111;
	assign font[13][9] = 14'b11111111111111;
	assign font[14][9] = 14'b11111111111111;
	assign font[15][9] = 14'b11111111111111;
	assign font[16][9] = 14'b11111111111111;
	assign font[17][9] = 14'b11111111111111;
	assign font[18][9] = 14'b11111111111111;
	assign font[19][9] = 14'b11111111111111;
	assign font[20][9] = 14'b11111111111111;
	assign font[21][9] = 14'b11111111111111;
	assign font[22][9] = 14'b11111111111111;
	assign font[23][9] = 14'b11111111111111;
	assign font[24][9] = 14'b11111111111111;
	assign font[25][9] = 14'b11111111111111;
	assign font[26][9] = 14'b11111111111111;
	assign font[27][9] = 14'b11111111111111;
	assign font[28][9] = 14'b11111111111111;
	assign font[29][9] = 14'b11111111111111;
	assign font[30][9] = 14'b11111111111111;
	assign font[31][9] = 14'b11111111111111;

	assign font[0][10] = 14'b11111111111111;
	assign font[1][10] = 14'b11111111111111;
	assign font[2][10] = 14'b11111111111111;
	assign font[3][10] = 14'b11111111111111;
	assign font[4][10] = 14'b11111111111111;
	assign font[5][10] = 14'b11111111111111;
	assign font[6][10] = 14'b11111111111111;
	assign font[7][10] = 14'b11111111111111;
	assign font[8][10] = 14'b11111111111111;
	assign font[9][10] = 14'b11111111111111;
	assign font[10][10] = 14'b11111111111111;
	assign font[11][10] = 14'b11111111111111;
	assign font[12][10] = 14'b11111111111111;
	assign font[13][10] = 14'b11111111111111;
	assign font[14][10] = 14'b11111111111111;
	assign font[15][10] = 14'b11111111111111;
	assign font[16][10] = 14'b11111111111111;
	assign font[17][10] = 14'b11111111111111;
	assign font[18][10] = 14'b11111111111111;
	assign font[19][10] = 14'b11111111111111;
	assign font[20][10] = 14'b11111111111111;
	assign font[21][10] = 14'b11111111111111;
	assign font[22][10] = 14'b11111111111111;
	assign font[23][10] = 14'b11111111111111;
	assign font[24][10] = 14'b11111111111111;
	assign font[25][10] = 14'b11111111111111;
	assign font[26][10] = 14'b11111111111111;
	assign font[27][10] = 14'b11111111111111;
	assign font[28][10] = 14'b11111111111111;
	assign font[29][10] = 14'b11111111111111;
	assign font[30][10] = 14'b11111111111111;
	assign font[31][10] = 14'b11111111111111;

	assign font[0][11] = 14'b11111111111111;
	assign font[1][11] = 14'b11111111111111;
	assign font[2][11] = 14'b11111111111111;
	assign font[3][11] = 14'b11111111111111;
	assign font[4][11] = 14'b11111111111111;
	assign font[5][11] = 14'b11111111111111;
	assign font[6][11] = 14'b11111111111111;
	assign font[7][11] = 14'b11111111111111;
	assign font[8][11] = 14'b11111111111111;
	assign font[9][11] = 14'b11111111111111;
	assign font[10][11] = 14'b11111111111111;
	assign font[11][11] = 14'b11111111111111;
	assign font[12][11] = 14'b11111111111111;
	assign font[13][11] = 14'b11111111111111;
	assign font[14][11] = 14'b11111111111111;
	assign font[15][11] = 14'b11111111111111;
	assign font[16][11] = 14'b11111111111111;
	assign font[17][11] = 14'b11111111111111;
	assign font[18][11] = 14'b11111111111111;
	assign font[19][11] = 14'b11111111111111;
	assign font[20][11] = 14'b11111111111111;
	assign font[21][11] = 14'b11111111111111;
	assign font[22][11] = 14'b11111111111111;
	assign font[23][11] = 14'b11111111111111;
	assign font[24][11] = 14'b11111111111111;
	assign font[25][11] = 14'b11111111111111;
	assign font[26][11] = 14'b11111111111111;
	assign font[27][11] = 14'b11111111111111;
	assign font[28][11] = 14'b11111111111111;
	assign font[29][11] = 14'b11111111111111;
	assign font[30][11] = 14'b11111111111111;
	assign font[31][11] = 14'b11111111111111;

	assign font[0][12] = 14'b11111111111111;
	assign font[1][12] = 14'b11111111111111;
	assign font[2][12] = 14'b11111111111111;
	assign font[3][12] = 14'b11111111111111;
	assign font[4][12] = 14'b11111111111111;
	assign font[5][12] = 14'b11111111111111;
	assign font[6][12] = 14'b11111111111111;
	assign font[7][12] = 14'b11111111111111;
	assign font[8][12] = 14'b11111111111111;
	assign font[9][12] = 14'b11111111111111;
	assign font[10][12] = 14'b11111111111111;
	assign font[11][12] = 14'b11111111111111;
	assign font[12][12] = 14'b11111111111111;
	assign font[13][12] = 14'b11111111111111;
	assign font[14][12] = 14'b11111111111111;
	assign font[15][12] = 14'b11111111111111;
	assign font[16][12] = 14'b11111111111111;
	assign font[17][12] = 14'b11111111111111;
	assign font[18][12] = 14'b11111111111111;
	assign font[19][12] = 14'b11111111111111;
	assign font[20][12] = 14'b11111111111111;
	assign font[21][12] = 14'b11111111111111;
	assign font[22][12] = 14'b11111111111111;
	assign font[23][12] = 14'b11111111111111;
	assign font[24][12] = 14'b11111111111111;
	assign font[25][12] = 14'b11111111111111;
	assign font[26][12] = 14'b11111111111111;
	assign font[27][12] = 14'b11111111111111;
	assign font[28][12] = 14'b11111111111111;
	assign font[29][12] = 14'b11111111111111;
	assign font[30][12] = 14'b11111111111111;
	assign font[31][12] = 14'b11111111111111;

	assign font[0][13] = 14'b11111111111111;
	assign font[1][13] = 14'b11111111111111;
	assign font[2][13] = 14'b11111111111111;
	assign font[3][13] = 14'b11111111111111;
	assign font[4][13] = 14'b11111111111111;
	assign font[5][13] = 14'b11111111111111;
	assign font[6][13] = 14'b11111111111111;
	assign font[7][13] = 14'b11111111111111;
	assign font[8][13] = 14'b11111111111111;
	assign font[9][13] = 14'b11111111111111;
	assign font[10][13] = 14'b11111111111111;
	assign font[11][13] = 14'b11111111111111;
	assign font[12][13] = 14'b11111111111111;
	assign font[13][13] = 14'b11111111111111;
	assign font[14][13] = 14'b11111111111111;
	assign font[15][13] = 14'b11111111111111;
	assign font[16][13] = 14'b11111111111111;
	assign font[17][13] = 14'b11111111111111;
	assign font[18][13] = 14'b11111111111111;
	assign font[19][13] = 14'b11111111111111;
	assign font[20][13] = 14'b11111111111111;
	assign font[21][13] = 14'b11111111111111;
	assign font[22][13] = 14'b11111111111111;
	assign font[23][13] = 14'b11111111111111;
	assign font[24][13] = 14'b11111111111111;
	assign font[25][13] = 14'b11111111111111;
	assign font[26][13] = 14'b11111111111111;
	assign font[27][13] = 14'b11111111111111;
	assign font[28][13] = 14'b11111111111111;
	assign font[29][13] = 14'b11111111111111;
	assign font[30][13] = 14'b11111111111111;
	assign font[31][13] = 14'b11111111111111;

	assign font[0][14] = 14'b11111111111111;
	assign font[1][14] = 14'b11111111111111;
	assign font[2][14] = 14'b11111111111111;
	assign font[3][14] = 14'b11111111111111;
	assign font[4][14] = 14'b11111111111111;
	assign font[5][14] = 14'b11111111111111;
	assign font[6][14] = 14'b11111111111111;
	assign font[7][14] = 14'b11111111111111;
	assign font[8][14] = 14'b11111111111111;
	assign font[9][14] = 14'b11111111111111;
	assign font[10][14] = 14'b11111111111111;
	assign font[11][14] = 14'b11111111111111;
	assign font[12][14] = 14'b11111111111111;
	assign font[13][14] = 14'b11111111111111;
	assign font[14][14] = 14'b11111111111111;
	assign font[15][14] = 14'b11111111111111;
	assign font[16][14] = 14'b11111111111111;
	assign font[17][14] = 14'b11111111111111;
	assign font[18][14] = 14'b11111111111111;
	assign font[19][14] = 14'b11111111111111;
	assign font[20][14] = 14'b11111111111111;
	assign font[21][14] = 14'b11111111111111;
	assign font[22][14] = 14'b11111111111111;
	assign font[23][14] = 14'b11111111111111;
	assign font[24][14] = 14'b11111111111111;
	assign font[25][14] = 14'b11111111111111;
	assign font[26][14] = 14'b11111111111111;
	assign font[27][14] = 14'b11111111111111;
	assign font[28][14] = 14'b11111111111111;
	assign font[29][14] = 14'b11111111111111;
	assign font[30][14] = 14'b11111111111111;
	assign font[31][14] = 14'b11111111111111;

	assign font[0][15] = 14'b11111111111111;
	assign font[1][15] = 14'b11111111111111;
	assign font[2][15] = 14'b11111111111111;
	assign font[3][15] = 14'b11111111111111;
	assign font[4][15] = 14'b11111111111111;
	assign font[5][15] = 14'b11111111111111;
	assign font[6][15] = 14'b11111111111111;
	assign font[7][15] = 14'b11111111111111;
	assign font[8][15] = 14'b11111111111111;
	assign font[9][15] = 14'b11111111111111;
	assign font[10][15] = 14'b11111111111111;
	assign font[11][15] = 14'b11111111111111;
	assign font[12][15] = 14'b11111111111111;
	assign font[13][15] = 14'b11111111111111;
	assign font[14][15] = 14'b11111111111111;
	assign font[15][15] = 14'b11111111111111;
	assign font[16][15] = 14'b11111111111111;
	assign font[17][15] = 14'b11111111111111;
	assign font[18][15] = 14'b11111111111111;
	assign font[19][15] = 14'b11111111111111;
	assign font[20][15] = 14'b11111111111111;
	assign font[21][15] = 14'b11111111111111;
	assign font[22][15] = 14'b11111111111111;
	assign font[23][15] = 14'b11111111111111;
	assign font[24][15] = 14'b11111111111111;
	assign font[25][15] = 14'b11111111111111;
	assign font[26][15] = 14'b11111111111111;
	assign font[27][15] = 14'b11111111111111;
	assign font[28][15] = 14'b11111111111111;
	assign font[29][15] = 14'b11111111111111;
	assign font[30][15] = 14'b11111111111111;
	assign font[31][15] = 14'b11111111111111;

	assign font[0][16] = 14'b11111111111111;
	assign font[1][16] = 14'b11111111111111;
	assign font[2][16] = 14'b11111111111111;
	assign font[3][16] = 14'b11111111111111;
	assign font[4][16] = 14'b11111111111111;
	assign font[5][16] = 14'b11111111111111;
	assign font[6][16] = 14'b11111111111111;
	assign font[7][16] = 14'b11111111111111;
	assign font[8][16] = 14'b11111111111111;
	assign font[9][16] = 14'b11111111111111;
	assign font[10][16] = 14'b11111111111111;
	assign font[11][16] = 14'b11111111111111;
	assign font[12][16] = 14'b11111111111111;
	assign font[13][16] = 14'b11111111111111;
	assign font[14][16] = 14'b11111111111111;
	assign font[15][16] = 14'b11111111111111;
	assign font[16][16] = 14'b11111111111111;
	assign font[17][16] = 14'b11111111111111;
	assign font[18][16] = 14'b11111111111111;
	assign font[19][16] = 14'b11111111111111;
	assign font[20][16] = 14'b11111111111111;
	assign font[21][16] = 14'b11111111111111;
	assign font[22][16] = 14'b11111111111111;
	assign font[23][16] = 14'b11111111111111;
	assign font[24][16] = 14'b11111111111111;
	assign font[25][16] = 14'b11111111111111;
	assign font[26][16] = 14'b11111111111111;
	assign font[27][16] = 14'b11111111111111;
	assign font[28][16] = 14'b11111111111111;
	assign font[29][16] = 14'b11111111111111;
	assign font[30][16] = 14'b11111111111111;
	assign font[31][16] = 14'b11111111111111;

	assign font[0][17] = 14'b11111111111111;
	assign font[1][17] = 14'b11111111111111;
	assign font[2][17] = 14'b11111111111111;
	assign font[3][17] = 14'b11111111111111;
	assign font[4][17] = 14'b11111111111111;
	assign font[5][17] = 14'b11111111111111;
	assign font[6][17] = 14'b11111111111111;
	assign font[7][17] = 14'b11111111111111;
	assign font[8][17] = 14'b11111111111111;
	assign font[9][17] = 14'b11111111111111;
	assign font[10][17] = 14'b11111111111111;
	assign font[11][17] = 14'b11111111111111;
	assign font[12][17] = 14'b11111111111111;
	assign font[13][17] = 14'b11111111111111;
	assign font[14][17] = 14'b11111111111111;
	assign font[15][17] = 14'b11111111111111;
	assign font[16][17] = 14'b11111111111111;
	assign font[17][17] = 14'b11111111111111;
	assign font[18][17] = 14'b11111111111111;
	assign font[19][17] = 14'b11111111111111;
	assign font[20][17] = 14'b11111111111111;
	assign font[21][17] = 14'b11111111111111;
	assign font[22][17] = 14'b11111111111111;
	assign font[23][17] = 14'b11111111111111;
	assign font[24][17] = 14'b11111111111111;
	assign font[25][17] = 14'b11111111111111;
	assign font[26][17] = 14'b11111111111111;
	assign font[27][17] = 14'b11111111111111;
	assign font[28][17] = 14'b11111111111111;
	assign font[29][17] = 14'b11111111111111;
	assign font[30][17] = 14'b11111111111111;
	assign font[31][17] = 14'b11111111111111;

	assign font[0][18] = 14'b11111111111111;
	assign font[1][18] = 14'b11111111111111;
	assign font[2][18] = 14'b11111111111111;
	assign font[3][18] = 14'b11111111111111;
	assign font[4][18] = 14'b11111111111111;
	assign font[5][18] = 14'b11111111111111;
	assign font[6][18] = 14'b11111111111111;
	assign font[7][18] = 14'b11111111111111;
	assign font[8][18] = 14'b11111111111111;
	assign font[9][18] = 14'b11111111111111;
	assign font[10][18] = 14'b11111111111111;
	assign font[11][18] = 14'b11111111111111;
	assign font[12][18] = 14'b11111111111111;
	assign font[13][18] = 14'b11111111111111;
	assign font[14][18] = 14'b11111111111111;
	assign font[15][18] = 14'b11111111111111;
	assign font[16][18] = 14'b11111111111111;
	assign font[17][18] = 14'b11111111111111;
	assign font[18][18] = 14'b11111111111111;
	assign font[19][18] = 14'b11111111111111;
	assign font[20][18] = 14'b11111111111111;
	assign font[21][18] = 14'b11111111111111;
	assign font[22][18] = 14'b11111111111111;
	assign font[23][18] = 14'b11111111111111;
	assign font[24][18] = 14'b11111111111111;
	assign font[25][18] = 14'b11111111111111;
	assign font[26][18] = 14'b11111111111111;
	assign font[27][18] = 14'b11111111111111;
	assign font[28][18] = 14'b11111111111111;
	assign font[29][18] = 14'b11111111111111;
	assign font[30][18] = 14'b11111111111111;
	assign font[31][18] = 14'b11111111111111;

	assign font[0][19] = 14'b11111111111111;
	assign font[1][19] = 14'b11111111111111;
	assign font[2][19] = 14'b11111111111111;
	assign font[3][19] = 14'b11111111111111;
	assign font[4][19] = 14'b11111111111111;
	assign font[5][19] = 14'b11111111111111;
	assign font[6][19] = 14'b11111111111111;
	assign font[7][19] = 14'b11111111111111;
	assign font[8][19] = 14'b11111111111111;
	assign font[9][19] = 14'b11111111111111;
	assign font[10][19] = 14'b11111111111111;
	assign font[11][19] = 14'b11111111111111;
	assign font[12][19] = 14'b11111111111111;
	assign font[13][19] = 14'b11111111111111;
	assign font[14][19] = 14'b11111111111111;
	assign font[15][19] = 14'b11111111111111;
	assign font[16][19] = 14'b11111111111111;
	assign font[17][19] = 14'b11111111111111;
	assign font[18][19] = 14'b11111111111111;
	assign font[19][19] = 14'b11111111111111;
	assign font[20][19] = 14'b11111111111111;
	assign font[21][19] = 14'b11111111111111;
	assign font[22][19] = 14'b11111111111111;
	assign font[23][19] = 14'b11111111111111;
	assign font[24][19] = 14'b11111111111111;
	assign font[25][19] = 14'b11111111111111;
	assign font[26][19] = 14'b11111111111111;
	assign font[27][19] = 14'b11111111111111;
	assign font[28][19] = 14'b11111111111111;
	assign font[29][19] = 14'b11111111111111;
	assign font[30][19] = 14'b11111111111111;
	assign font[31][19] = 14'b11111111111111;

	assign font[0][20] = 14'b11111111111111;
	assign font[1][20] = 14'b11111111111111;
	assign font[2][20] = 14'b11111111111111;
	assign font[3][20] = 14'b11111111111111;
	assign font[4][20] = 14'b11111111111111;
	assign font[5][20] = 14'b11111111111111;
	assign font[6][20] = 14'b11111111111111;
	assign font[7][20] = 14'b11111111111111;
	assign font[8][20] = 14'b11111111111111;
	assign font[9][20] = 14'b11111111111111;
	assign font[10][20] = 14'b11111111111111;
	assign font[11][20] = 14'b11111111111111;
	assign font[12][20] = 14'b11111111111111;
	assign font[13][20] = 14'b11111111111111;
	assign font[14][20] = 14'b11111111111111;
	assign font[15][20] = 14'b11111111111111;
	assign font[16][20] = 14'b11111111111111;
	assign font[17][20] = 14'b11111111111111;
	assign font[18][20] = 14'b11111111111111;
	assign font[19][20] = 14'b11111111111111;
	assign font[20][20] = 14'b11111111111111;
	assign font[21][20] = 14'b11111111111111;
	assign font[22][20] = 14'b11111111111111;
	assign font[23][20] = 14'b11111111111111;
	assign font[24][20] = 14'b11111111111111;
	assign font[25][20] = 14'b11111111111111;
	assign font[26][20] = 14'b11111111111111;
	assign font[27][20] = 14'b11111111111111;
	assign font[28][20] = 14'b11111111111111;
	assign font[29][20] = 14'b11111111111111;
	assign font[30][20] = 14'b11111111111111;
	assign font[31][20] = 14'b11111111111111;

	assign font[0][21] = 14'b11111111111111;
	assign font[1][21] = 14'b11111111111111;
	assign font[2][21] = 14'b11111111111111;
	assign font[3][21] = 14'b11111111111111;
	assign font[4][21] = 14'b11111111111111;
	assign font[5][21] = 14'b11111111111111;
	assign font[6][21] = 14'b11111111111111;
	assign font[7][21] = 14'b11111111111111;
	assign font[8][21] = 14'b11111111111111;
	assign font[9][21] = 14'b11111111111111;
	assign font[10][21] = 14'b11111111111111;
	assign font[11][21] = 14'b11111111111111;
	assign font[12][21] = 14'b11111111111111;
	assign font[13][21] = 14'b11111111111111;
	assign font[14][21] = 14'b11111111111111;
	assign font[15][21] = 14'b11111111111111;
	assign font[16][21] = 14'b11111111111111;
	assign font[17][21] = 14'b11111111111111;
	assign font[18][21] = 14'b11111111111111;
	assign font[19][21] = 14'b11111111111111;
	assign font[20][21] = 14'b11111111111111;
	assign font[21][21] = 14'b11111111111111;
	assign font[22][21] = 14'b11111111111111;
	assign font[23][21] = 14'b11111111111111;
	assign font[24][21] = 14'b11111111111111;
	assign font[25][21] = 14'b11111111111111;
	assign font[26][21] = 14'b11111111111111;
	assign font[27][21] = 14'b11111111111111;
	assign font[28][21] = 14'b11111111111111;
	assign font[29][21] = 14'b11111111111111;
	assign font[30][21] = 14'b11111111111111;
	assign font[31][21] = 14'b11111111111111;

	assign font[0][22] = 14'b11111111111111;
	assign font[1][22] = 14'b11111111111111;
	assign font[2][22] = 14'b11111111111111;
	assign font[3][22] = 14'b11111111111111;
	assign font[4][22] = 14'b11111111111111;
	assign font[5][22] = 14'b11111111111111;
	assign font[6][22] = 14'b11111111111111;
	assign font[7][22] = 14'b11111111111111;
	assign font[8][22] = 14'b11111111111111;
	assign font[9][22] = 14'b11111111111111;
	assign font[10][22] = 14'b11111111111111;
	assign font[11][22] = 14'b11111111111111;
	assign font[12][22] = 14'b11111111111111;
	assign font[13][22] = 14'b11111111111111;
	assign font[14][22] = 14'b11111111111111;
	assign font[15][22] = 14'b11111111111111;
	assign font[16][22] = 14'b11111111111111;
	assign font[17][22] = 14'b11111111111111;
	assign font[18][22] = 14'b11111111111111;
	assign font[19][22] = 14'b11111111111111;
	assign font[20][22] = 14'b11111111111111;
	assign font[21][22] = 14'b11111111111111;
	assign font[22][22] = 14'b11111111111111;
	assign font[23][22] = 14'b11111111111111;
	assign font[24][22] = 14'b11111111111111;
	assign font[25][22] = 14'b11111111111111;
	assign font[26][22] = 14'b11111111111111;
	assign font[27][22] = 14'b11111111111111;
	assign font[28][22] = 14'b11111111111111;
	assign font[29][22] = 14'b11111111111111;
	assign font[30][22] = 14'b11111111111111;
	assign font[31][22] = 14'b11111111111111;

	assign font[0][23] = 14'b11111111111111;
	assign font[1][23] = 14'b11111111111111;
	assign font[2][23] = 14'b11111111111111;
	assign font[3][23] = 14'b11111111111111;
	assign font[4][23] = 14'b11111111111111;
	assign font[5][23] = 14'b11111111111111;
	assign font[6][23] = 14'b11111111111111;
	assign font[7][23] = 14'b11111111111111;
	assign font[8][23] = 14'b11111111111111;
	assign font[9][23] = 14'b11111111111111;
	assign font[10][23] = 14'b11111111111111;
	assign font[11][23] = 14'b11111111111111;
	assign font[12][23] = 14'b11111111111111;
	assign font[13][23] = 14'b11111111111111;
	assign font[14][23] = 14'b11111111111111;
	assign font[15][23] = 14'b11111111111111;
	assign font[16][23] = 14'b11111111111111;
	assign font[17][23] = 14'b11111111111111;
	assign font[18][23] = 14'b11111111111111;
	assign font[19][23] = 14'b11111111111111;
	assign font[20][23] = 14'b11111111111111;
	assign font[21][23] = 14'b11111111111111;
	assign font[22][23] = 14'b11111111111111;
	assign font[23][23] = 14'b11111111111111;
	assign font[24][23] = 14'b11111111111111;
	assign font[25][23] = 14'b11111111111111;
	assign font[26][23] = 14'b11111111111111;
	assign font[27][23] = 14'b11111111111111;
	assign font[28][23] = 14'b11111111111111;
	assign font[29][23] = 14'b11111111111111;
	assign font[30][23] = 14'b11111111111111;
	assign font[31][23] = 14'b11111111111111;

	assign font[0][24] = 14'b11111111111111;
	assign font[1][24] = 14'b11111111111111;
	assign font[2][24] = 14'b11111111111111;
	assign font[3][24] = 14'b11111111111111;
	assign font[4][24] = 14'b11111111111111;
	assign font[5][24] = 14'b11111111111111;
	assign font[6][24] = 14'b11111111111111;
	assign font[7][24] = 14'b11111111111111;
	assign font[8][24] = 14'b11111111111111;
	assign font[9][24] = 14'b11111111111111;
	assign font[10][24] = 14'b11111111111111;
	assign font[11][24] = 14'b11111111111111;
	assign font[12][24] = 14'b11111111111111;
	assign font[13][24] = 14'b11111111111111;
	assign font[14][24] = 14'b11111111111111;
	assign font[15][24] = 14'b11111111111111;
	assign font[16][24] = 14'b11111111111111;
	assign font[17][24] = 14'b11111111111111;
	assign font[18][24] = 14'b11111111111111;
	assign font[19][24] = 14'b11111111111111;
	assign font[20][24] = 14'b11111111111111;
	assign font[21][24] = 14'b11111111111111;
	assign font[22][24] = 14'b11111111111111;
	assign font[23][24] = 14'b11111111111111;
	assign font[24][24] = 14'b11111111111111;
	assign font[25][24] = 14'b11111111111111;
	assign font[26][24] = 14'b11111111111111;
	assign font[27][24] = 14'b11111111111111;
	assign font[28][24] = 14'b11111111111111;
	assign font[29][24] = 14'b11111111111111;
	assign font[30][24] = 14'b11111111111111;
	assign font[31][24] = 14'b11111111111111;

	assign font[0][25] = 14'b11111111111111;
	assign font[1][25] = 14'b11111111111111;
	assign font[2][25] = 14'b11111111111111;
	assign font[3][25] = 14'b11111111111111;
	assign font[4][25] = 14'b11111111111111;
	assign font[5][25] = 14'b11111111111111;
	assign font[6][25] = 14'b11111111111111;
	assign font[7][25] = 14'b11111111111111;
	assign font[8][25] = 14'b11111111111111;
	assign font[9][25] = 14'b11111111111111;
	assign font[10][25] = 14'b11111111111111;
	assign font[11][25] = 14'b11111111111111;
	assign font[12][25] = 14'b11111111111111;
	assign font[13][25] = 14'b11111111111111;
	assign font[14][25] = 14'b11111111111111;
	assign font[15][25] = 14'b11111111111111;
	assign font[16][25] = 14'b11111111111111;
	assign font[17][25] = 14'b11111111111111;
	assign font[18][25] = 14'b11111111111111;
	assign font[19][25] = 14'b11111111111111;
	assign font[20][25] = 14'b11111111111111;
	assign font[21][25] = 14'b11111111111111;
	assign font[22][25] = 14'b11111111111111;
	assign font[23][25] = 14'b11111111111111;
	assign font[24][25] = 14'b11111111111111;
	assign font[25][25] = 14'b11111111111111;
	assign font[26][25] = 14'b11111111111111;
	assign font[27][25] = 14'b11111111111111;
	assign font[28][25] = 14'b11111111111111;
	assign font[29][25] = 14'b11111111111111;
	assign font[30][25] = 14'b11111111111111;
	assign font[31][25] = 14'b11111111111111;

	assign font[0][26] = 14'b11111111111111;
	assign font[1][26] = 14'b11111111111111;
	assign font[2][26] = 14'b11111111111111;
	assign font[3][26] = 14'b11111111111111;
	assign font[4][26] = 14'b11111111111111;
	assign font[5][26] = 14'b11111111111111;
	assign font[6][26] = 14'b11111111111111;
	assign font[7][26] = 14'b11111111111111;
	assign font[8][26] = 14'b11111111111111;
	assign font[9][26] = 14'b11111111111111;
	assign font[10][26] = 14'b11111111111111;
	assign font[11][26] = 14'b11111111111111;
	assign font[12][26] = 14'b11111111111111;
	assign font[13][26] = 14'b11111111111111;
	assign font[14][26] = 14'b11111111111111;
	assign font[15][26] = 14'b11111111111111;
	assign font[16][26] = 14'b11111111111111;
	assign font[17][26] = 14'b11111111111111;
	assign font[18][26] = 14'b11111111111111;
	assign font[19][26] = 14'b11111111111111;
	assign font[20][26] = 14'b11111111111111;
	assign font[21][26] = 14'b11111111111111;
	assign font[22][26] = 14'b11111111111111;
	assign font[23][26] = 14'b11111111111111;
	assign font[24][26] = 14'b11111111111111;
	assign font[25][26] = 14'b11111111111111;
	assign font[26][26] = 14'b11111111111111;
	assign font[27][26] = 14'b11111111111111;
	assign font[28][26] = 14'b11111111111111;
	assign font[29][26] = 14'b11111111111111;
	assign font[30][26] = 14'b11111111111111;
	assign font[31][26] = 14'b11111111111111;

	assign font[0][27] = 14'b11111111111111;
	assign font[1][27] = 14'b11111111111111;
	assign font[2][27] = 14'b11111111111111;
	assign font[3][27] = 14'b11111111111111;
	assign font[4][27] = 14'b11111111111111;
	assign font[5][27] = 14'b11111111111111;
	assign font[6][27] = 14'b11111111111111;
	assign font[7][27] = 14'b11111111111111;
	assign font[8][27] = 14'b11111111111111;
	assign font[9][27] = 14'b11111111111111;
	assign font[10][27] = 14'b11111111111111;
	assign font[11][27] = 14'b11111111111111;
	assign font[12][27] = 14'b11111111111111;
	assign font[13][27] = 14'b11111111111111;
	assign font[14][27] = 14'b11111111111111;
	assign font[15][27] = 14'b11111111111111;
	assign font[16][27] = 14'b11111111111111;
	assign font[17][27] = 14'b11111111111111;
	assign font[18][27] = 14'b11111111111111;
	assign font[19][27] = 14'b11111111111111;
	assign font[20][27] = 14'b11111111111111;
	assign font[21][27] = 14'b11111111111111;
	assign font[22][27] = 14'b11111111111111;
	assign font[23][27] = 14'b11111111111111;
	assign font[24][27] = 14'b11111111111111;
	assign font[25][27] = 14'b11111111111111;
	assign font[26][27] = 14'b11111111111111;
	assign font[27][27] = 14'b11111111111111;
	assign font[28][27] = 14'b11111111111111;
	assign font[29][27] = 14'b11111111111111;
	assign font[30][27] = 14'b11111111111111;
	assign font[31][27] = 14'b11111111111111;

	assign font[0][28] = 14'b11111111111111;
	assign font[1][28] = 14'b11111111111111;
	assign font[2][28] = 14'b11111111111111;
	assign font[3][28] = 14'b11111111111111;
	assign font[4][28] = 14'b11111111111111;
	assign font[5][28] = 14'b11111111111111;
	assign font[6][28] = 14'b11111111111111;
	assign font[7][28] = 14'b11111111111111;
	assign font[8][28] = 14'b11111111111111;
	assign font[9][28] = 14'b11111111111111;
	assign font[10][28] = 14'b11111111111111;
	assign font[11][28] = 14'b11111111111111;
	assign font[12][28] = 14'b11111111111111;
	assign font[13][28] = 14'b11111111111111;
	assign font[14][28] = 14'b11111111111111;
	assign font[15][28] = 14'b11111111111111;
	assign font[16][28] = 14'b11111111111111;
	assign font[17][28] = 14'b11111111111111;
	assign font[18][28] = 14'b11111111111111;
	assign font[19][28] = 14'b11111111111111;
	assign font[20][28] = 14'b11111111111111;
	assign font[21][28] = 14'b11111111111111;
	assign font[22][28] = 14'b11111111111111;
	assign font[23][28] = 14'b11111111111111;
	assign font[24][28] = 14'b11111111111111;
	assign font[25][28] = 14'b11111111111111;
	assign font[26][28] = 14'b11111111111111;
	assign font[27][28] = 14'b11111111111111;
	assign font[28][28] = 14'b11111111111111;
	assign font[29][28] = 14'b11111111111111;
	assign font[30][28] = 14'b11111111111111;
	assign font[31][28] = 14'b11111111111111;

	assign font[0][29] = 14'b11111111111111;
	assign font[1][29] = 14'b11111111111111;
	assign font[2][29] = 14'b11111111111111;
	assign font[3][29] = 14'b11111111111111;
	assign font[4][29] = 14'b11111111111111;
	assign font[5][29] = 14'b11111111111111;
	assign font[6][29] = 14'b11111111111111;
	assign font[7][29] = 14'b11111111111111;
	assign font[8][29] = 14'b11111111111111;
	assign font[9][29] = 14'b11111111111111;
	assign font[10][29] = 14'b11111111111111;
	assign font[11][29] = 14'b11111111111111;
	assign font[12][29] = 14'b11111111111111;
	assign font[13][29] = 14'b11111111111111;
	assign font[14][29] = 14'b11111111111111;
	assign font[15][29] = 14'b11111111111111;
	assign font[16][29] = 14'b11111111111111;
	assign font[17][29] = 14'b11111111111111;
	assign font[18][29] = 14'b11111111111111;
	assign font[19][29] = 14'b11111111111111;
	assign font[20][29] = 14'b11111111111111;
	assign font[21][29] = 14'b11111111111111;
	assign font[22][29] = 14'b11111111111111;
	assign font[23][29] = 14'b11111111111111;
	assign font[24][29] = 14'b11111111111111;
	assign font[25][29] = 14'b11111111111111;
	assign font[26][29] = 14'b11111111111111;
	assign font[27][29] = 14'b11111111111111;
	assign font[28][29] = 14'b11111111111111;
	assign font[29][29] = 14'b11111111111111;
	assign font[30][29] = 14'b11111111111111;
	assign font[31][29] = 14'b11111111111111;

	assign font[0][30] = 14'b11111111111111;
	assign font[1][30] = 14'b11111111111111;
	assign font[2][30] = 14'b11111111111111;
	assign font[3][30] = 14'b11111111111111;
	assign font[4][30] = 14'b11111111111111;
	assign font[5][30] = 14'b11111111111111;
	assign font[6][30] = 14'b11111111111111;
	assign font[7][30] = 14'b11111111111111;
	assign font[8][30] = 14'b11111111111111;
	assign font[9][30] = 14'b11111111111111;
	assign font[10][30] = 14'b11111111111111;
	assign font[11][30] = 14'b11111111111111;
	assign font[12][30] = 14'b11111111111111;
	assign font[13][30] = 14'b11111111111111;
	assign font[14][30] = 14'b11111111111111;
	assign font[15][30] = 14'b11111111111111;
	assign font[16][30] = 14'b11111111111111;
	assign font[17][30] = 14'b11111111111111;
	assign font[18][30] = 14'b11111111111111;
	assign font[19][30] = 14'b11111111111111;
	assign font[20][30] = 14'b11111111111111;
	assign font[21][30] = 14'b11111111111111;
	assign font[22][30] = 14'b11111111111111;
	assign font[23][30] = 14'b11111111111111;
	assign font[24][30] = 14'b11111111111111;
	assign font[25][30] = 14'b11111111111111;
	assign font[26][30] = 14'b11111111111111;
	assign font[27][30] = 14'b11111111111111;
	assign font[28][30] = 14'b11111111111111;
	assign font[29][30] = 14'b11111111111111;
	assign font[30][30] = 14'b11111111111111;
	assign font[31][30] = 14'b11111111111111;

	assign font[0][31] = 14'b11111111111111;
	assign font[1][31] = 14'b11111111111111;
	assign font[2][31] = 14'b11111111111111;
	assign font[3][31] = 14'b11111111111111;
	assign font[4][31] = 14'b11111111111111;
	assign font[5][31] = 14'b11111111111111;
	assign font[6][31] = 14'b11111111111111;
	assign font[7][31] = 14'b11111111111111;
	assign font[8][31] = 14'b11111111111111;
	assign font[9][31] = 14'b11111111111111;
	assign font[10][31] = 14'b11111111111111;
	assign font[11][31] = 14'b11111111111111;
	assign font[12][31] = 14'b11111111111111;
	assign font[13][31] = 14'b11111111111111;
	assign font[14][31] = 14'b11111111111111;
	assign font[15][31] = 14'b11111111111111;
	assign font[16][31] = 14'b11111111111111;
	assign font[17][31] = 14'b11111111111111;
	assign font[18][31] = 14'b11111111111111;
	assign font[19][31] = 14'b11111111111111;
	assign font[20][31] = 14'b11111111111111;
	assign font[21][31] = 14'b11111111111111;
	assign font[22][31] = 14'b11111111111111;
	assign font[23][31] = 14'b11111111111111;
	assign font[24][31] = 14'b11111111111111;
	assign font[25][31] = 14'b11111111111111;
	assign font[26][31] = 14'b11111111111111;
	assign font[27][31] = 14'b11111111111111;
	assign font[28][31] = 14'b11111111111111;
	assign font[29][31] = 14'b11111111111111;
	assign font[30][31] = 14'b11111111111111;
	assign font[31][31] = 14'b11111111111111;

	assign font[0][32] = 14'b11111111111111;
	assign font[1][32] = 14'b11111111111111;
	assign font[2][32] = 14'b11111111111111;
	assign font[3][32] = 14'b11111111111111;
	assign font[4][32] = 14'b11111111111111;
	assign font[5][32] = 14'b11111111111111;
	assign font[6][32] = 14'b11111111111111;
	assign font[7][32] = 14'b11111111111111;
	assign font[8][32] = 14'b11111111111111;
	assign font[9][32] = 14'b11111111111111;
	assign font[10][32] = 14'b11111111111111;
	assign font[11][32] = 14'b11111111111111;
	assign font[12][32] = 14'b11111111111111;
	assign font[13][32] = 14'b11111111111111;
	assign font[14][32] = 14'b11111111111111;
	assign font[15][32] = 14'b11111111111111;
	assign font[16][32] = 14'b11111111111111;
	assign font[17][32] = 14'b11111111111111;
	assign font[18][32] = 14'b11111111111111;
	assign font[19][32] = 14'b11111111111111;
	assign font[20][32] = 14'b11111111111111;
	assign font[21][32] = 14'b11111111111111;
	assign font[22][32] = 14'b11111111111111;
	assign font[23][32] = 14'b11111111111111;
	assign font[24][32] = 14'b11111111111111;
	assign font[25][32] = 14'b11111111111111;
	assign font[26][32] = 14'b11111111111111;
	assign font[27][32] = 14'b11111111111111;
	assign font[28][32] = 14'b11111111111111;
	assign font[29][32] = 14'b11111111111111;
	assign font[30][32] = 14'b11111111111111;
	assign font[31][32] = 14'b11111111111111;

	assign font[0][33] = 14'b00000000000000;
	assign font[1][33] = 14'b00000000000000;
	assign font[2][33] = 14'b00000000000000;
	assign font[3][33] = 14'b00000000000000;
	assign font[4][33] = 14'b00000000000000;
	assign font[5][33] = 14'b00000000000000;
	assign font[6][33] = 14'b00000000000000;
	assign font[7][33] = 14'b00000000000000;
	assign font[8][33] = 14'b00000000000000;
	assign font[9][33] = 14'b00000011100000;
	assign font[10][33] = 14'b00000011100000;
	assign font[11][33] = 14'b00000011100000;
	assign font[12][33] = 14'b00000011100000;
	assign font[13][33] = 14'b00000011100000;
	assign font[14][33] = 14'b00000011100000;
	assign font[15][33] = 14'b00000011100000;
	assign font[16][33] = 14'b00000011100000;
	assign font[17][33] = 14'b00000011100000;
	assign font[18][33] = 14'b00000011100000;
	assign font[19][33] = 14'b00000011100000;
	assign font[20][33] = 14'b00000011100000;
	assign font[21][33] = 14'b00000011100000;
	assign font[22][33] = 14'b00000000000000;
	assign font[23][33] = 14'b00000000000000;
	assign font[24][33] = 14'b00000000000000;
	assign font[25][33] = 14'b00000011100000;
	assign font[26][33] = 14'b00000011100000;
	assign font[27][33] = 14'b00000000000000;
	assign font[28][33] = 14'b00000000000000;
	assign font[29][33] = 14'b00000000000000;
	assign font[30][33] = 14'b00000000000000;
	assign font[31][33] = 14'b00000000000000;

	assign font[0][34] = 14'b00000000000000;
	assign font[1][34] = 14'b00000000000000;
	assign font[2][34] = 14'b00000000000000;
	assign font[3][34] = 14'b00000000000000;
	assign font[4][34] = 14'b00000000000000;
	assign font[5][34] = 14'b00000000000000;
	assign font[6][34] = 14'b00011100111000;
	assign font[7][34] = 14'b00011100111000;
	assign font[8][34] = 14'b00011100111000;
	assign font[9][34] = 14'b00011100111000;
	assign font[10][34] = 14'b00011100111000;
	assign font[11][34] = 14'b00000000000000;
	assign font[12][34] = 14'b00000000000000;
	assign font[13][34] = 14'b00000000000000;
	assign font[14][34] = 14'b00000000000000;
	assign font[15][34] = 14'b00000000000000;
	assign font[16][34] = 14'b00000000000000;
	assign font[17][34] = 14'b00000000000000;
	assign font[18][34] = 14'b00000000000000;
	assign font[19][34] = 14'b00000000000000;
	assign font[20][34] = 14'b00000000000000;
	assign font[21][34] = 14'b00000000000000;
	assign font[22][34] = 14'b00000000000000;
	assign font[23][34] = 14'b00000000000000;
	assign font[24][34] = 14'b00000000000000;
	assign font[25][34] = 14'b00000000000000;
	assign font[26][34] = 14'b00000000000000;
	assign font[27][34] = 14'b00000000000000;
	assign font[28][34] = 14'b00000000000000;
	assign font[29][34] = 14'b00000000000000;
	assign font[30][34] = 14'b00000000000000;
	assign font[31][34] = 14'b00000000000000;

	assign font[0][35] = 14'b00000000000000;
	assign font[1][35] = 14'b00000000000000;
	assign font[2][35] = 14'b00000000000000;
	assign font[3][35] = 14'b00000000000000;
	assign font[4][35] = 14'b00000000000000;
	assign font[5][35] = 14'b00000000000000;
	assign font[6][35] = 14'b00000000000000;
	assign font[7][35] = 14'b00000000000000;
	assign font[8][35] = 14'b00000000000000;
	assign font[9][35] = 14'b00000000000000;
	assign font[10][35] = 14'b00000000000000;
	assign font[11][35] = 14'b00000000000000;
	assign font[12][35] = 14'b00001110111000;
	assign font[13][35] = 14'b00001110111000;
	assign font[14][35] = 14'b00111111111110;
	assign font[15][35] = 14'b00111111111110;
	assign font[16][35] = 14'b00001110111000;
	assign font[17][35] = 14'b00001110111000;
	assign font[18][35] = 14'b00001110111000;
	assign font[19][35] = 14'b00001110111000;
	assign font[20][35] = 14'b00001110111000;
	assign font[21][35] = 14'b00001110111000;
	assign font[22][35] = 14'b00111111111110;
	assign font[23][35] = 14'b00111111111110;
	assign font[24][35] = 14'b00001110111000;
	assign font[25][35] = 14'b00001110111000;
	assign font[26][35] = 14'b00001110111000;
	assign font[27][35] = 14'b00000000000000;
	assign font[28][35] = 14'b00000000000000;
	assign font[29][35] = 14'b00000000000000;
	assign font[30][35] = 14'b00000000000000;
	assign font[31][35] = 14'b00000000000000;

	assign font[0][36] = 14'b00000000000000;
	assign font[1][36] = 14'b00000000000000;
	assign font[2][36] = 14'b00000000000000;
	assign font[3][36] = 14'b00000000000000;
	assign font[4][36] = 14'b00000000000000;
	assign font[5][36] = 14'b00000000000000;
	assign font[6][36] = 14'b00000000000000;
	assign font[7][36] = 14'b00000000000000;
	assign font[8][36] = 14'b00000000000000;
	assign font[9][36] = 14'b00000011000000;
	assign font[10][36] = 14'b00000011000000;
	assign font[11][36] = 14'b00000011000000;
	assign font[12][36] = 14'b00001111111000;
	assign font[13][36] = 14'b00001111111000;
	assign font[14][36] = 14'b00111011000000;
	assign font[15][36] = 14'b00111011000000;
	assign font[16][36] = 14'b00001111111000;
	assign font[17][36] = 14'b00001111111000;
	assign font[18][36] = 14'b00001111111000;
	assign font[19][36] = 14'b00000011001110;
	assign font[20][36] = 14'b00000011001110;
	assign font[21][36] = 14'b00000011001000;
	assign font[22][36] = 14'b00001111111000;
	assign font[23][36] = 14'b00001111111000;
	assign font[24][36] = 14'b00000011000000;
	assign font[25][36] = 14'b00000011000000;
	assign font[26][36] = 14'b00000011000000;
	assign font[27][36] = 14'b00000000000000;
	assign font[28][36] = 14'b00000000000000;
	assign font[29][36] = 14'b00000000000000;
	assign font[30][36] = 14'b00000000000000;
	assign font[31][36] = 14'b00000000000000;

	assign font[0][37] = 14'b00000000000000;
	assign font[1][37] = 14'b00000000000000;
	assign font[2][37] = 14'b00000000000000;
	assign font[3][37] = 14'b00000000000000;
	assign font[4][37] = 14'b00000000000000;
	assign font[5][37] = 14'b00000000000000;
	assign font[6][37] = 14'b00000000000000;
	assign font[7][37] = 14'b00000000000000;
	assign font[8][37] = 14'b00000000000000;
	assign font[9][37] = 14'b00011100011000;
	assign font[10][37] = 14'b00011100011000;
	assign font[11][37] = 14'b00010100010000;
	assign font[12][37] = 14'b00110110110000;
	assign font[13][37] = 14'b00110110110000;
	assign font[14][37] = 14'b00011100100000;
	assign font[15][37] = 14'b00011101100000;
	assign font[16][37] = 14'b00011100100000;
	assign font[17][37] = 14'b00000001000000;
	assign font[18][37] = 14'b00000001100000;
	assign font[19][37] = 14'b00000011011100;
	assign font[20][37] = 14'b00000011011100;
	assign font[21][37] = 14'b00000011011100;
	assign font[22][37] = 14'b00000110110110;
	assign font[23][37] = 14'b00000110110110;
	assign font[24][37] = 14'b00000100010100;
	assign font[25][37] = 14'b00001100011100;
	assign font[26][37] = 14'b00001100011100;
	assign font[27][37] = 14'b00000000000000;
	assign font[28][37] = 14'b00000000000000;
	assign font[29][37] = 14'b00000000000000;
	assign font[30][37] = 14'b00000000000000;
	assign font[31][37] = 14'b00000000000000;

	assign font[0][38] = 14'b00000000000000;
	assign font[1][38] = 14'b00000000000000;
	assign font[2][38] = 14'b00000000000000;
	assign font[3][38] = 14'b00000000000000;
	assign font[4][38] = 14'b00000000000000;
	assign font[5][38] = 14'b00000000000000;
	assign font[6][38] = 14'b00000000000000;
	assign font[7][38] = 14'b00000000000000;
	assign font[8][38] = 14'b00000000000000;
	assign font[9][38] = 14'b00000111100000;
	assign font[10][38] = 14'b00000111100000;
	assign font[11][38] = 14'b00001100110000;
	assign font[12][38] = 14'b00001100110000;
	assign font[13][38] = 14'b00001100110000;
	assign font[14][38] = 14'b00000111100110;
	assign font[15][38] = 14'b00000111100110;
	assign font[16][38] = 14'b00011111100110;
	assign font[17][38] = 14'b00011101100110;
	assign font[18][38] = 14'b00011101100110;
	assign font[19][38] = 14'b00111000111000;
	assign font[20][38] = 14'b00111000111000;
	assign font[21][38] = 14'b00111000111100;
	assign font[22][38] = 14'b00111001101100;
	assign font[23][38] = 14'b00111001101100;
	assign font[24][38] = 14'b00001001101100;
	assign font[25][38] = 14'b00001111101110;
	assign font[26][38] = 14'b00001111101110;
	assign font[27][38] = 14'b00000000000000;
	assign font[28][38] = 14'b00000000000000;
	assign font[29][38] = 14'b00000000000000;
	assign font[30][38] = 14'b00000000000000;
	assign font[31][38] = 14'b00000000000000;

	assign font[0][39] = 14'b00000000000000;
	assign font[1][39] = 14'b00000000000000;
	assign font[2][39] = 14'b00000000000000;
	assign font[3][39] = 14'b00000000000000;
	assign font[4][39] = 14'b00000000000000;
	assign font[5][39] = 14'b00000000000000;
	assign font[6][39] = 14'b00000000000000;
	assign font[7][39] = 14'b00000011100000;
	assign font[8][39] = 14'b00000011100000;
	assign font[9][39] = 14'b00001110000000;
	assign font[10][39] = 14'b00001110000000;
	assign font[11][39] = 14'b00001110000000;
	assign font[12][39] = 14'b00000000000000;
	assign font[13][39] = 14'b00000000000000;
	assign font[14][39] = 14'b00000000000000;
	assign font[15][39] = 14'b00000000000000;
	assign font[16][39] = 14'b00000000000000;
	assign font[17][39] = 14'b00000000000000;
	assign font[18][39] = 14'b00000000000000;
	assign font[19][39] = 14'b00000000000000;
	assign font[20][39] = 14'b00000000000000;
	assign font[21][39] = 14'b00000000000000;
	assign font[22][39] = 14'b00000000000000;
	assign font[23][39] = 14'b00000000000000;
	assign font[24][39] = 14'b00000000000000;
	assign font[25][39] = 14'b00000000000000;
	assign font[26][39] = 14'b00000000000000;
	assign font[27][39] = 14'b00000000000000;
	assign font[28][39] = 14'b00000000000000;
	assign font[29][39] = 14'b00000000000000;
	assign font[30][39] = 14'b00000000000000;
	assign font[31][39] = 14'b00000000000000;

	assign font[0][40] = 14'b00000000000000;
	assign font[1][40] = 14'b00000000000000;
	assign font[2][40] = 14'b00000000000000;
	assign font[3][40] = 14'b00000000000000;
	assign font[4][40] = 14'b00000000000000;
	assign font[5][40] = 14'b00000000000000;
	assign font[6][40] = 14'b00000000110000;
	assign font[7][40] = 14'b00000000110000;
	assign font[8][40] = 14'b00000000000000;
	assign font[9][40] = 14'b00000011000000;
	assign font[10][40] = 14'b00000011000000;
	assign font[11][40] = 14'b00000110000000;
	assign font[12][40] = 14'b00000110000000;
	assign font[13][40] = 14'b00000110000000;
	assign font[14][40] = 14'b00001110000000;
	assign font[15][40] = 14'b00001110000000;
	assign font[16][40] = 14'b00001110000000;
	assign font[17][40] = 14'b00001110000000;
	assign font[18][40] = 14'b00001110000000;
	assign font[19][40] = 14'b00001110000000;
	assign font[20][40] = 14'b00001110000000;
	assign font[21][40] = 14'b00001110000000;
	assign font[22][40] = 14'b00000110000000;
	assign font[23][40] = 14'b00000110000000;
	assign font[24][40] = 14'b00000011000000;
	assign font[25][40] = 14'b00000011000000;
	assign font[26][40] = 14'b00000011000000;
	assign font[27][40] = 14'b00000000110000;
	assign font[28][40] = 14'b00000000110000;
	assign font[29][40] = 14'b00000000000000;
	assign font[30][40] = 14'b00000000000000;
	assign font[31][40] = 14'b00000000000000;

	assign font[0][41] = 14'b00000000000000;
	assign font[1][41] = 14'b00000000000000;
	assign font[2][41] = 14'b00000000000000;
	assign font[3][41] = 14'b00000000000000;
	assign font[4][41] = 14'b00000000000000;
	assign font[5][41] = 14'b00000000000000;
	assign font[6][41] = 14'b00001100000000;
	assign font[7][41] = 14'b00001100000000;
	assign font[8][41] = 14'b00000000000000;
	assign font[9][41] = 14'b00000011000000;
	assign font[10][41] = 14'b00000011000000;
	assign font[11][41] = 14'b00000001100000;
	assign font[12][41] = 14'b00000001100000;
	assign font[13][41] = 14'b00000001100000;
	assign font[14][41] = 14'b00000001110000;
	assign font[15][41] = 14'b00000001110000;
	assign font[16][41] = 14'b00000001110000;
	assign font[17][41] = 14'b00000001110000;
	assign font[18][41] = 14'b00000001110000;
	assign font[19][41] = 14'b00000001110000;
	assign font[20][41] = 14'b00000001110000;
	assign font[21][41] = 14'b00000001110000;
	assign font[22][41] = 14'b00000001100000;
	assign font[23][41] = 14'b00000001100000;
	assign font[24][41] = 14'b00000001000000;
	assign font[25][41] = 14'b00000011000000;
	assign font[26][41] = 14'b00000011000000;
	assign font[27][41] = 14'b00001100000000;
	assign font[28][41] = 14'b00001100000000;
	assign font[29][41] = 14'b00001100000000;
	assign font[30][41] = 14'b00000000000000;
	assign font[31][41] = 14'b00000000000000;

	assign font[0][42] = 14'b00000000000000;
	assign font[1][42] = 14'b00000000000000;
	assign font[2][42] = 14'b00000000000000;
	assign font[3][42] = 14'b00000000000000;
	assign font[4][42] = 14'b00000000000000;
	assign font[5][42] = 14'b00000000000000;
	assign font[6][42] = 14'b00000000000000;
	assign font[7][42] = 14'b00000000000000;
	assign font[8][42] = 14'b00000000000000;
	assign font[9][42] = 14'b00000000000000;
	assign font[10][42] = 14'b00000000000000;
	assign font[11][42] = 14'b00000010000000;
	assign font[12][42] = 14'b00000011000000;
	assign font[13][42] = 14'b00000011000000;
	assign font[14][42] = 14'b00111011111000;
	assign font[15][42] = 14'b00111011111000;
	assign font[16][42] = 14'b00000011000000;
	assign font[17][42] = 14'b00000111000000;
	assign font[18][42] = 14'b00000111000000;
	assign font[19][42] = 14'b00111011111000;
	assign font[20][42] = 14'b00111011111000;
	assign font[21][42] = 14'b00111011111000;
	assign font[22][42] = 14'b00000011000000;
	assign font[23][42] = 14'b00000011000000;
	assign font[24][42] = 14'b00000011000000;
	assign font[25][42] = 14'b00000000000000;
	assign font[26][42] = 14'b00000000000000;
	assign font[27][42] = 14'b00000000000000;
	assign font[28][42] = 14'b00000000000000;
	assign font[29][42] = 14'b00000000000000;
	assign font[30][42] = 14'b00000000000000;
	assign font[31][42] = 14'b00000000000000;

	assign font[0][43] = 14'b00000000000000;
	assign font[1][43] = 14'b00000000000000;
	assign font[2][43] = 14'b00000000000000;
	assign font[3][43] = 14'b00000000000000;
	assign font[4][43] = 14'b00000000000000;
	assign font[5][43] = 14'b00000000000000;
	assign font[6][43] = 14'b00000000000000;
	assign font[7][43] = 14'b00000000000000;
	assign font[8][43] = 14'b00000000000000;
	assign font[9][43] = 14'b00000000000000;
	assign font[10][43] = 14'b00000000000000;
	assign font[11][43] = 14'b00000011100000;
	assign font[12][43] = 14'b00000011100000;
	assign font[13][43] = 14'b00000011100000;
	assign font[14][43] = 14'b00000011100000;
	assign font[15][43] = 14'b00000011100000;
	assign font[16][43] = 14'b00111111111100;
	assign font[17][43] = 14'b00011111111100;
	assign font[18][43] = 14'b00000011100000;
	assign font[19][43] = 14'b00000011100000;
	assign font[20][43] = 14'b00000011100000;
	assign font[21][43] = 14'b00000011100000;
	assign font[22][43] = 14'b00000011100000;
	assign font[23][43] = 14'b00000011100000;
	assign font[24][43] = 14'b00000000000000;
	assign font[25][43] = 14'b00000000000000;
	assign font[26][43] = 14'b00000000000000;
	assign font[27][43] = 14'b00000000000000;
	assign font[28][43] = 14'b00000000000000;
	assign font[29][43] = 14'b00000000000000;
	assign font[30][43] = 14'b00000000000000;
	assign font[31][43] = 14'b00000000000000;

	assign font[0][44] = 14'b00000000000000;
	assign font[1][44] = 14'b00000000000000;
	assign font[2][44] = 14'b00000000000000;
	assign font[3][44] = 14'b00000000000000;
	assign font[4][44] = 14'b00000000000000;
	assign font[5][44] = 14'b00000000000000;
	assign font[6][44] = 14'b00000000000000;
	assign font[7][44] = 14'b00000000000000;
	assign font[8][44] = 14'b00000000000000;
	assign font[9][44] = 14'b00000000000000;
	assign font[10][44] = 14'b00000000000000;
	assign font[11][44] = 14'b00000000000000;
	assign font[12][44] = 14'b00000000000000;
	assign font[13][44] = 14'b00000000000000;
	assign font[14][44] = 14'b00000000000000;
	assign font[15][44] = 14'b00000000000000;
	assign font[16][44] = 14'b00000000000000;
	assign font[17][44] = 14'b00000000000000;
	assign font[18][44] = 14'b00000000000000;
	assign font[19][44] = 14'b00000000000000;
	assign font[20][44] = 14'b00000000000000;
	assign font[21][44] = 14'b00000000000000;
	assign font[22][44] = 14'b00000011110000;
	assign font[23][44] = 14'b00000011110000;
	assign font[24][44] = 14'b00000011110000;
	assign font[25][44] = 14'b00000011110000;
	assign font[26][44] = 14'b00000011110000;
	assign font[27][44] = 14'b00000111100000;
	assign font[28][44] = 14'b00000111100000;
	assign font[29][44] = 14'b00000111100000;
	assign font[30][44] = 14'b00011110000000;
	assign font[31][44] = 14'b00011110000000;

	assign font[0][45] = 14'b00000000000000;
	assign font[1][45] = 14'b00000000000000;
	assign font[2][45] = 14'b00000000000000;
	assign font[3][45] = 14'b00000000000000;
	assign font[4][45] = 14'b00000000000000;
	assign font[5][45] = 14'b00000000000000;
	assign font[6][45] = 14'b00000000000000;
	assign font[7][45] = 14'b00000000000000;
	assign font[8][45] = 14'b00000000000000;
	assign font[9][45] = 14'b00000000000000;
	assign font[10][45] = 14'b00000000000000;
	assign font[11][45] = 14'b00000000000000;
	assign font[12][45] = 14'b00000000000000;
	assign font[13][45] = 14'b00000000000000;
	assign font[14][45] = 14'b00000000000000;
	assign font[15][45] = 14'b00000000000000;
	assign font[16][45] = 14'b00000000000000;
	assign font[17][45] = 14'b00011111111000;
	assign font[18][45] = 14'b00011111111000;
	assign font[19][45] = 14'b00000000000000;
	assign font[20][45] = 14'b00000000000000;
	assign font[21][45] = 14'b00000000000000;
	assign font[22][45] = 14'b00000000000000;
	assign font[23][45] = 14'b00000000000000;
	assign font[24][45] = 14'b00000000000000;
	assign font[25][45] = 14'b00000000000000;
	assign font[26][45] = 14'b00000000000000;
	assign font[27][45] = 14'b00000000000000;
	assign font[28][45] = 14'b00000000000000;
	assign font[29][45] = 14'b00000000000000;
	assign font[30][45] = 14'b00000000000000;
	assign font[31][45] = 14'b00000000000000;

	assign font[0][46] = 14'b00000000000000;
	assign font[1][46] = 14'b00000000000000;
	assign font[2][46] = 14'b00000000000000;
	assign font[3][46] = 14'b00000000000000;
	assign font[4][46] = 14'b00000000000000;
	assign font[5][46] = 14'b00000000000000;
	assign font[6][46] = 14'b00000000000000;
	assign font[7][46] = 14'b00000000000000;
	assign font[8][46] = 14'b00000000000000;
	assign font[9][46] = 14'b00000000000000;
	assign font[10][46] = 14'b00000000000000;
	assign font[11][46] = 14'b00000000000000;
	assign font[12][46] = 14'b00000000000000;
	assign font[13][46] = 14'b00000000000000;
	assign font[14][46] = 14'b00000000000000;
	assign font[15][46] = 14'b00000000000000;
	assign font[16][46] = 14'b00000000000000;
	assign font[17][46] = 14'b00000000000000;
	assign font[18][46] = 14'b00000000000000;
	assign font[19][46] = 14'b00000000000000;
	assign font[20][46] = 14'b00000000000000;
	assign font[21][46] = 14'b00000000000000;
	assign font[22][46] = 14'b00000111100000;
	assign font[23][46] = 14'b00000111100000;
	assign font[24][46] = 14'b00000111100000;
	assign font[25][46] = 14'b00000111100000;
	assign font[26][46] = 14'b00000111100000;
	assign font[27][46] = 14'b00000000000000;
	assign font[28][46] = 14'b00000000000000;
	assign font[29][46] = 14'b00000000000000;
	assign font[30][46] = 14'b00000000000000;
	assign font[31][46] = 14'b00000000000000;

	assign font[0][47] = 14'b00000000000000;
	assign font[1][47] = 14'b00000000000000;
	assign font[2][47] = 14'b00000000000000;
	assign font[3][47] = 14'b00000000000000;
	assign font[4][47] = 14'b00000000000000;
	assign font[5][47] = 14'b00000000000000;
	assign font[6][47] = 14'b00000000001110;
	assign font[7][47] = 14'b00000000001110;
	assign font[8][47] = 14'b00000000001110;
	assign font[9][47] = 14'b00000000011100;
	assign font[10][47] = 14'b00000000011100;
	assign font[11][47] = 14'b00000000111000;
	assign font[12][47] = 14'b00000000111000;
	assign font[13][47] = 14'b00000000111000;
	assign font[14][47] = 14'b00000001110000;
	assign font[15][47] = 14'b00000001110000;
	assign font[16][47] = 14'b00000001110000;
	assign font[17][47] = 14'b00000001100000;
	assign font[18][47] = 14'b00000001100000;
	assign font[19][47] = 14'b00000011100000;
	assign font[20][47] = 14'b00000011100000;
	assign font[21][47] = 14'b00000011100000;
	assign font[22][47] = 14'b00000111000000;
	assign font[23][47] = 14'b00000111000000;
	assign font[24][47] = 14'b00000110000000;
	assign font[25][47] = 14'b00001110000000;
	assign font[26][47] = 14'b00001110000000;
	assign font[27][47] = 14'b00011100000000;
	assign font[28][47] = 14'b00011100000000;
	assign font[29][47] = 14'b00000000000000;
	assign font[30][47] = 14'b00000000000000;
	assign font[31][47] = 14'b00000000000000;

	assign font[0][48] = 14'b00000000000000;
	assign font[1][48] = 14'b00000000000000;
	assign font[2][48] = 14'b00000000000000;
	assign font[3][48] = 14'b00000000000000;
	assign font[4][48] = 14'b00000000000000;
	assign font[5][48] = 14'b00000000000000;
	assign font[6][48] = 14'b00000000000000;
	assign font[7][48] = 14'b00000000000000;
	assign font[8][48] = 14'b00000000000000;
	assign font[9][48] = 14'b00000011110000;
	assign font[10][48] = 14'b00000011110000;
	assign font[11][48] = 14'b00001100011000;
	assign font[12][48] = 14'b00001100011000;
	assign font[13][48] = 14'b00001100011000;
	assign font[14][48] = 14'b00011100011100;
	assign font[15][48] = 14'b00011100011100;
	assign font[16][48] = 14'b00011100011100;
	assign font[17][48] = 14'b00011100011100;
	assign font[18][48] = 14'b00011100011100;
	assign font[19][48] = 14'b00011100011100;
	assign font[20][48] = 14'b00011100011100;
	assign font[21][48] = 14'b00011100011100;
	assign font[22][48] = 14'b00001100011000;
	assign font[23][48] = 14'b00001100011000;
	assign font[24][48] = 14'b00000000000000;
	assign font[25][48] = 14'b00000011110000;
	assign font[26][48] = 14'b00000011110000;
	assign font[27][48] = 14'b00000000000000;
	assign font[28][48] = 14'b00000000000000;
	assign font[29][48] = 14'b00000000000000;
	assign font[30][48] = 14'b00000000000000;
	assign font[31][48] = 14'b00000000000000;

	assign font[0][49] = 14'b00000000000000;
	assign font[1][49] = 14'b00000000000000;
	assign font[2][49] = 14'b00000000000000;
	assign font[3][49] = 14'b00000000000000;
	assign font[4][49] = 14'b00000000000000;
	assign font[5][49] = 14'b00000000000000;
	assign font[6][49] = 14'b00000000000000;
	assign font[7][49] = 14'b00000000000000;
	assign font[8][49] = 14'b00000000000000;
	assign font[9][49] = 14'b00000011100000;
	assign font[10][49] = 14'b00000011100000;
	assign font[11][49] = 14'b00000011100000;
	assign font[12][49] = 14'b00001111100000;
	assign font[13][49] = 14'b00001111100000;
	assign font[14][49] = 14'b00000011100000;
	assign font[15][49] = 14'b00000011100000;
	assign font[16][49] = 14'b00000011100000;
	assign font[17][49] = 14'b00000011100000;
	assign font[18][49] = 14'b00000011100000;
	assign font[19][49] = 14'b00000011100000;
	assign font[20][49] = 14'b00000011100000;
	assign font[21][49] = 14'b00000011100000;
	assign font[22][49] = 14'b00000011100000;
	assign font[23][49] = 14'b00000011100000;
	assign font[24][49] = 14'b00000011100000;
	assign font[25][49] = 14'b00011111111000;
	assign font[26][49] = 14'b00011111111000;
	assign font[27][49] = 14'b00000000000000;
	assign font[28][49] = 14'b00000000000000;
	assign font[29][49] = 14'b00000000000000;
	assign font[30][49] = 14'b00000000000000;
	assign font[31][49] = 14'b00000000000000;

	assign font[0][50] = 14'b00000000000000;
	assign font[1][50] = 14'b00000000000000;
	assign font[2][50] = 14'b00000000000000;
	assign font[3][50] = 14'b00000000000000;
	assign font[4][50] = 14'b00000000000000;
	assign font[5][50] = 14'b00000000000000;
	assign font[6][50] = 14'b00000000000000;
	assign font[7][50] = 14'b00000000000000;
	assign font[8][50] = 14'b00000000000000;
	assign font[9][50] = 14'b00001111110000;
	assign font[10][50] = 14'b00001111110000;
	assign font[11][50] = 14'b00011000011100;
	assign font[12][50] = 14'b00011000011100;
	assign font[13][50] = 14'b00000000011100;
	assign font[14][50] = 14'b00000000011100;
	assign font[15][50] = 14'b00000000011100;
	assign font[16][50] = 14'b00000000111000;
	assign font[17][50] = 14'b00000000111000;
	assign font[18][50] = 14'b00000000111000;
	assign font[19][50] = 14'b00000001110000;
	assign font[20][50] = 14'b00000001110000;
	assign font[21][50] = 14'b00000001110000;
	assign font[22][50] = 14'b00000111000000;
	assign font[23][50] = 14'b00000111000000;
	assign font[24][50] = 14'b00000111000000;
	assign font[25][50] = 14'b00011111111100;
	assign font[26][50] = 14'b00011111111100;
	assign font[27][50] = 14'b00000000000000;
	assign font[28][50] = 14'b00000000000000;
	assign font[29][50] = 14'b00000000000000;
	assign font[30][50] = 14'b00000000000000;
	assign font[31][50] = 14'b00000000000000;

	assign font[0][51] = 14'b00000000000000;
	assign font[1][51] = 14'b00000000000000;
	assign font[2][51] = 14'b00000000000000;
	assign font[3][51] = 14'b00000000000000;
	assign font[4][51] = 14'b00000000000000;
	assign font[5][51] = 14'b00000000000000;
	assign font[6][51] = 14'b00000000000000;
	assign font[7][51] = 14'b00000000000000;
	assign font[8][51] = 14'b00000000000000;
	assign font[9][51] = 14'b00001111110000;
	assign font[10][51] = 14'b00001111110000;
	assign font[11][51] = 14'b00111000011100;
	assign font[12][51] = 14'b00111000011100;
	assign font[13][51] = 14'b00000000011100;
	assign font[14][51] = 14'b00000000011100;
	assign font[15][51] = 14'b00000000011100;
	assign font[16][51] = 14'b00000000010000;
	assign font[17][51] = 14'b00000111110000;
	assign font[18][51] = 14'b00000111110000;
	assign font[19][51] = 14'b00000000011100;
	assign font[20][51] = 14'b00000000011100;
	assign font[21][51] = 14'b00000000011100;
	assign font[22][51] = 14'b00111000011100;
	assign font[23][51] = 14'b00111000011100;
	assign font[24][51] = 14'b00001000010000;
	assign font[25][51] = 14'b00001111110000;
	assign font[26][51] = 14'b00001111110000;
	assign font[27][51] = 14'b00000000000000;
	assign font[28][51] = 14'b00000000000000;
	assign font[29][51] = 14'b00000000000000;
	assign font[30][51] = 14'b00000000000000;
	assign font[31][51] = 14'b00000000000000;

	assign font[0][52] = 14'b00000000000000;
	assign font[1][52] = 14'b00000000000000;
	assign font[2][52] = 14'b00000000000000;
	assign font[3][52] = 14'b00000000000000;
	assign font[4][52] = 14'b00000000000000;
	assign font[5][52] = 14'b00000000000000;
	assign font[6][52] = 14'b00000000000000;
	assign font[7][52] = 14'b00000000000000;
	assign font[8][52] = 14'b00000000000000;
	assign font[9][52] = 14'b00000011110000;
	assign font[10][52] = 14'b00000011110000;
	assign font[11][52] = 14'b00000001110000;
	assign font[12][52] = 14'b00001101110000;
	assign font[13][52] = 14'b00001101110000;
	assign font[14][52] = 14'b00011001110000;
	assign font[15][52] = 14'b00011001110000;
	assign font[16][52] = 14'b00011001110000;
	assign font[17][52] = 14'b00110001110000;
	assign font[18][52] = 14'b00110001110000;
	assign font[19][52] = 14'b01111111111100;
	assign font[20][52] = 14'b01111111111100;
	assign font[21][52] = 14'b00000001110000;
	assign font[22][52] = 14'b00000001110000;
	assign font[23][52] = 14'b00000001110000;
	assign font[24][52] = 14'b00000001110000;
	assign font[25][52] = 14'b00000001110000;
	assign font[26][52] = 14'b00000001110000;
	assign font[27][52] = 14'b00000000000000;
	assign font[28][52] = 14'b00000000000000;
	assign font[29][52] = 14'b00000000000000;
	assign font[30][52] = 14'b00000000000000;
	assign font[31][52] = 14'b00000000000000;

	assign font[0][53] = 14'b00000000000000;
	assign font[1][53] = 14'b00000000000000;
	assign font[2][53] = 14'b00000000000000;
	assign font[3][53] = 14'b00000000000000;
	assign font[4][53] = 14'b00000000000000;
	assign font[5][53] = 14'b00000000000000;
	assign font[6][53] = 14'b00000000000000;
	assign font[7][53] = 14'b00000000000000;
	assign font[8][53] = 14'b00000000000000;
	assign font[9][53] = 14'b00111111111000;
	assign font[10][53] = 14'b00111111111000;
	assign font[11][53] = 14'b00111000000000;
	assign font[12][53] = 14'b00111000000000;
	assign font[13][53] = 14'b00111000000000;
	assign font[14][53] = 14'b00111011110000;
	assign font[15][53] = 14'b00111011110000;
	assign font[16][53] = 14'b00111100111000;
	assign font[17][53] = 14'b00111100111000;
	assign font[18][53] = 14'b00111100111000;
	assign font[19][53] = 14'b00000000011100;
	assign font[20][53] = 14'b00000000011100;
	assign font[21][53] = 14'b00000000011100;
	assign font[22][53] = 14'b00110000111000;
	assign font[23][53] = 14'b00110000111000;
	assign font[24][53] = 14'b00000000110000;
	assign font[25][53] = 14'b00001111110000;
	assign font[26][53] = 14'b00001111110000;
	assign font[27][53] = 14'b00000000000000;
	assign font[28][53] = 14'b00000000000000;
	assign font[29][53] = 14'b00000000000000;
	assign font[30][53] = 14'b00000000000000;
	assign font[31][53] = 14'b00000000000000;

	assign font[0][54] = 14'b00000000000000;
	assign font[1][54] = 14'b00000000000000;
	assign font[2][54] = 14'b00000000000000;
	assign font[3][54] = 14'b00000000000000;
	assign font[4][54] = 14'b00000000000000;
	assign font[5][54] = 14'b00000000000000;
	assign font[6][54] = 14'b00000000000000;
	assign font[7][54] = 14'b00000000000000;
	assign font[8][54] = 14'b00000000000000;
	assign font[9][54] = 14'b00000011111000;
	assign font[10][54] = 14'b00000011111000;
	assign font[11][54] = 14'b00000000000000;
	assign font[12][54] = 14'b00001110000000;
	assign font[13][54] = 14'b00001110000000;
	assign font[14][54] = 14'b00011100000000;
	assign font[15][54] = 14'b00011100000000;
	assign font[16][54] = 14'b00011100000000;
	assign font[17][54] = 14'b00011111111000;
	assign font[18][54] = 14'b00011111111000;
	assign font[19][54] = 14'b00011110001110;
	assign font[20][54] = 14'b00011110001110;
	assign font[21][54] = 14'b00001110001110;
	assign font[22][54] = 14'b00001110001110;
	assign font[23][54] = 14'b00001110001110;
	assign font[24][54] = 14'b00000000001000;
	assign font[25][54] = 14'b00000011111000;
	assign font[26][54] = 14'b00000011111000;
	assign font[27][54] = 14'b00000000000000;
	assign font[28][54] = 14'b00000000000000;
	assign font[29][54] = 14'b00000000000000;
	assign font[30][54] = 14'b00000000000000;
	assign font[31][54] = 14'b00000000000000;

	assign font[0][55] = 14'b00000000000000;
	assign font[1][55] = 14'b00000000000000;
	assign font[2][55] = 14'b00000000000000;
	assign font[3][55] = 14'b00000000000000;
	assign font[4][55] = 14'b00000000000000;
	assign font[5][55] = 14'b00000000000000;
	assign font[6][55] = 14'b00000000000000;
	assign font[7][55] = 14'b00000000000000;
	assign font[8][55] = 14'b00000000000000;
	assign font[9][55] = 14'b00111111111000;
	assign font[10][55] = 14'b00111111111000;
	assign font[11][55] = 14'b00000000111000;
	assign font[12][55] = 14'b00000000111000;
	assign font[13][55] = 14'b00000000111000;
	assign font[14][55] = 14'b00000001110000;
	assign font[15][55] = 14'b00000001110000;
	assign font[16][55] = 14'b00000001110000;
	assign font[17][55] = 14'b00000011100000;
	assign font[18][55] = 14'b00000011100000;
	assign font[19][55] = 14'b00000011000000;
	assign font[20][55] = 14'b00000111000000;
	assign font[21][55] = 14'b00000111000000;
	assign font[22][55] = 14'b00000110000000;
	assign font[23][55] = 14'b00000110000000;
	assign font[24][55] = 14'b00001110000000;
	assign font[25][55] = 14'b00001110000000;
	assign font[26][55] = 14'b00001110000000;
	assign font[27][55] = 14'b00000000000000;
	assign font[28][55] = 14'b00000000000000;
	assign font[29][55] = 14'b00000000000000;
	assign font[30][55] = 14'b00000000000000;
	assign font[31][55] = 14'b00000000000000;

	assign font[0][56] = 14'b00000000000000;
	assign font[1][56] = 14'b00000000000000;
	assign font[2][56] = 14'b00000000000000;
	assign font[3][56] = 14'b00000000000000;
	assign font[4][56] = 14'b00000000000000;
	assign font[5][56] = 14'b00000000000000;
	assign font[6][56] = 14'b00000000000000;
	assign font[7][56] = 14'b00000000000000;
	assign font[8][56] = 14'b00000000000000;
	assign font[9][56] = 14'b00000111111000;
	assign font[10][56] = 14'b00000111111000;
	assign font[11][56] = 14'b00011100011100;
	assign font[12][56] = 14'b00011100011100;
	assign font[13][56] = 14'b00011100011100;
	assign font[14][56] = 14'b00011100011100;
	assign font[15][56] = 14'b00011100011100;
	assign font[16][56] = 14'b00001100011000;
	assign font[17][56] = 14'b00001111111000;
	assign font[18][56] = 14'b00001111111000;
	assign font[19][56] = 14'b00011100011100;
	assign font[20][56] = 14'b00011100011100;
	assign font[21][56] = 14'b00011100011100;
	assign font[22][56] = 14'b00011100011100;
	assign font[23][56] = 14'b00011100011100;
	assign font[24][56] = 14'b00000100011000;
	assign font[25][56] = 14'b00000111111000;
	assign font[26][56] = 14'b00000111111000;
	assign font[27][56] = 14'b00000000000000;
	assign font[28][56] = 14'b00000000000000;
	assign font[29][56] = 14'b00000000000000;
	assign font[30][56] = 14'b00000000000000;
	assign font[31][56] = 14'b00000000000000;

	assign font[0][57] = 14'b00000000000000;
	assign font[1][57] = 14'b00000000000000;
	assign font[2][57] = 14'b00000000000000;
	assign font[3][57] = 14'b00000000000000;
	assign font[4][57] = 14'b00000000000000;
	assign font[5][57] = 14'b00000000000000;
	assign font[6][57] = 14'b00000000000000;
	assign font[7][57] = 14'b00000000000000;
	assign font[8][57] = 14'b00000000000000;
	assign font[9][57] = 14'b00001111110000;
	assign font[10][57] = 14'b00001111110000;
	assign font[11][57] = 14'b00111000111000;
	assign font[12][57] = 14'b00111000111000;
	assign font[13][57] = 14'b00111000111000;
	assign font[14][57] = 14'b00111000111100;
	assign font[15][57] = 14'b00111000111100;
	assign font[16][57] = 14'b00111000111100;
	assign font[17][57] = 14'b00001111111100;
	assign font[18][57] = 14'b00001111111100;
	assign font[19][57] = 14'b00000000011100;
	assign font[20][57] = 14'b00000000011100;
	assign font[21][57] = 14'b00000000011100;
	assign font[22][57] = 14'b00000000111000;
	assign font[23][57] = 14'b00000000111000;
	assign font[24][57] = 14'b00000000110000;
	assign font[25][57] = 14'b00001111110000;
	assign font[26][57] = 14'b00001111110000;
	assign font[27][57] = 14'b00000000000000;
	assign font[28][57] = 14'b00000000000000;
	assign font[29][57] = 14'b00000000000000;
	assign font[30][57] = 14'b00000000000000;
	assign font[31][57] = 14'b00000000000000;

	assign font[0][58] = 14'b00000000000000;
	assign font[1][58] = 14'b00000000000000;
	assign font[2][58] = 14'b00000000000000;
	assign font[3][58] = 14'b00000000000000;
	assign font[4][58] = 14'b00000000000000;
	assign font[5][58] = 14'b00000000000000;
	assign font[6][58] = 14'b00000000000000;
	assign font[7][58] = 14'b00000000000000;
	assign font[8][58] = 14'b00000000000000;
	assign font[9][58] = 14'b00000000000000;
	assign font[10][58] = 14'b00000000000000;
	assign font[11][58] = 14'b00000111100000;
	assign font[12][58] = 14'b00000111100000;
	assign font[13][58] = 14'b00000111100000;
	assign font[14][58] = 14'b00000111100000;
	assign font[15][58] = 14'b00000111100000;
	assign font[16][58] = 14'b00000000000000;
	assign font[17][58] = 14'b00000000000000;
	assign font[18][58] = 14'b00000000000000;
	assign font[19][58] = 14'b00000000000000;
	assign font[20][58] = 14'b00000000000000;
	assign font[21][58] = 14'b00000000000000;
	assign font[22][58] = 14'b00000111100000;
	assign font[23][58] = 14'b00000111100000;
	assign font[24][58] = 14'b00000111100000;
	assign font[25][58] = 14'b00000111100000;
	assign font[26][58] = 14'b00000111100000;
	assign font[27][58] = 14'b00000000000000;
	assign font[28][58] = 14'b00000000000000;
	assign font[29][58] = 14'b00000000000000;
	assign font[30][58] = 14'b00000000000000;
	assign font[31][58] = 14'b00000000000000;

	assign font[0][59] = 14'b00000000000000;
	assign font[1][59] = 14'b00000000000000;
	assign font[2][59] = 14'b00000000000000;
	assign font[3][59] = 14'b00000000000000;
	assign font[4][59] = 14'b00000000000000;
	assign font[5][59] = 14'b00000000000000;
	assign font[6][59] = 14'b00000000000000;
	assign font[7][59] = 14'b00000000000000;
	assign font[8][59] = 14'b00000000000000;
	assign font[9][59] = 14'b00000000000000;
	assign font[10][59] = 14'b00000000000000;
	assign font[11][59] = 14'b00000111100000;
	assign font[12][59] = 14'b00000111100000;
	assign font[13][59] = 14'b00000111100000;
	assign font[14][59] = 14'b00000111100000;
	assign font[15][59] = 14'b00000111100000;
	assign font[16][59] = 14'b00000000000000;
	assign font[17][59] = 14'b00000000000000;
	assign font[18][59] = 14'b00000000000000;
	assign font[19][59] = 14'b00000000000000;
	assign font[20][59] = 14'b00000000000000;
	assign font[21][59] = 14'b00000000000000;
	assign font[22][59] = 14'b00000111100000;
	assign font[23][59] = 14'b00000111100000;
	assign font[24][59] = 14'b00000111100000;
	assign font[25][59] = 14'b00000111100000;
	assign font[26][59] = 14'b00000111100000;
	assign font[27][59] = 14'b00001111000000;
	assign font[28][59] = 14'b00001111000000;
	assign font[29][59] = 14'b00001111000000;
	assign font[30][59] = 14'b00111100000000;
	assign font[31][59] = 14'b00111100000000;

	assign font[0][60] = 14'b00000000000000;
	assign font[1][60] = 14'b00000000000000;
	assign font[2][60] = 14'b00000000000000;
	assign font[3][60] = 14'b00000000000000;
	assign font[4][60] = 14'b00000000000000;
	assign font[5][60] = 14'b00000000000000;
	assign font[6][60] = 14'b00000000000000;
	assign font[7][60] = 14'b00000000000000;
	assign font[8][60] = 14'b00000000000000;
	assign font[9][60] = 14'b00000000111000;
	assign font[10][60] = 14'b00000000111000;
	assign font[11][60] = 14'b00000001110000;
	assign font[12][60] = 14'b00000001110000;
	assign font[13][60] = 14'b00000001110000;
	assign font[14][60] = 14'b00000111000000;
	assign font[15][60] = 14'b00000111000000;
	assign font[16][60] = 14'b00011100000000;
	assign font[17][60] = 14'b00011100000000;
	assign font[18][60] = 14'b00011100000000;
	assign font[19][60] = 14'b00000111000000;
	assign font[20][60] = 14'b00000111000000;
	assign font[21][60] = 14'b00000111000000;
	assign font[22][60] = 14'b00000001110000;
	assign font[23][60] = 14'b00000001110000;
	assign font[24][60] = 14'b00000000110000;
	assign font[25][60] = 14'b00000000111000;
	assign font[26][60] = 14'b00000000111000;
	assign font[27][60] = 14'b00000000000000;
	assign font[28][60] = 14'b00000000000000;
	assign font[29][60] = 14'b00000000000000;
	assign font[30][60] = 14'b00000000000000;
	assign font[31][60] = 14'b00000000000000;

	assign font[0][61] = 14'b00000000000000;
	assign font[1][61] = 14'b00000000000000;
	assign font[2][61] = 14'b00000000000000;
	assign font[3][61] = 14'b00000000000000;
	assign font[4][61] = 14'b00000000000000;
	assign font[5][61] = 14'b00000000000000;
	assign font[6][61] = 14'b00000000000000;
	assign font[7][61] = 14'b00000000000000;
	assign font[8][61] = 14'b00000000000000;
	assign font[9][61] = 14'b00000000000000;
	assign font[10][61] = 14'b00000000000000;
	assign font[11][61] = 14'b00000000000000;
	assign font[12][61] = 14'b00000000000000;
	assign font[13][61] = 14'b00000000000000;
	assign font[14][61] = 14'b00011111111000;
	assign font[15][61] = 14'b00011111111000;
	assign font[16][61] = 14'b00000000000000;
	assign font[17][61] = 14'b00000000000000;
	assign font[18][61] = 14'b00000000000000;
	assign font[19][61] = 14'b00011111111000;
	assign font[20][61] = 14'b00011111111000;
	assign font[21][61] = 14'b00000000000000;
	assign font[22][61] = 14'b00000000000000;
	assign font[23][61] = 14'b00000000000000;
	assign font[24][61] = 14'b00000000000000;
	assign font[25][61] = 14'b00000000000000;
	assign font[26][61] = 14'b00000000000000;
	assign font[27][61] = 14'b00000000000000;
	assign font[28][61] = 14'b00000000000000;
	assign font[29][61] = 14'b00000000000000;
	assign font[30][61] = 14'b00000000000000;
	assign font[31][61] = 14'b00000000000000;

	assign font[0][62] = 14'b00000000000000;
	assign font[1][62] = 14'b00000000000000;
	assign font[2][62] = 14'b00000000000000;
	assign font[3][62] = 14'b00000000000000;
	assign font[4][62] = 14'b00000000000000;
	assign font[5][62] = 14'b00000000000000;
	assign font[6][62] = 14'b00000000000000;
	assign font[7][62] = 14'b00000000000000;
	assign font[8][62] = 14'b00000000000000;
	assign font[9][62] = 14'b00111000000000;
	assign font[10][62] = 14'b00111000000000;
	assign font[11][62] = 14'b00001110000000;
	assign font[12][62] = 14'b00001110000000;
	assign font[13][62] = 14'b00001110000000;
	assign font[14][62] = 14'b00000011100000;
	assign font[15][62] = 14'b00000011100000;
	assign font[16][62] = 14'b00000001100000;
	assign font[17][62] = 14'b00000001110000;
	assign font[18][62] = 14'b00000001110000;
	assign font[19][62] = 14'b00000011100000;
	assign font[20][62] = 14'b00000011100000;
	assign font[21][62] = 14'b00000011100000;
	assign font[22][62] = 14'b00001110000000;
	assign font[23][62] = 14'b00001110000000;
	assign font[24][62] = 14'b00001000000000;
	assign font[25][62] = 14'b00111000000000;
	assign font[26][62] = 14'b00111000000000;
	assign font[27][62] = 14'b00000000000000;
	assign font[28][62] = 14'b00000000000000;
	assign font[29][62] = 14'b00000000000000;
	assign font[30][62] = 14'b00000000000000;
	assign font[31][62] = 14'b00000000000000;

	assign font[0][63] = 14'b00000000000000;
	assign font[1][63] = 14'b00000000000000;
	assign font[2][63] = 14'b00000000000000;
	assign font[3][63] = 14'b00000000000000;
	assign font[4][63] = 14'b00000000000000;
	assign font[5][63] = 14'b00000000000000;
	assign font[6][63] = 14'b00000000000000;
	assign font[7][63] = 14'b00000000000000;
	assign font[8][63] = 14'b00000000000000;
	assign font[9][63] = 14'b00001111110000;
	assign font[10][63] = 14'b00001111110000;
	assign font[11][63] = 14'b00001000110000;
	assign font[12][63] = 14'b00111000111000;
	assign font[13][63] = 14'b00111000111000;
	assign font[14][63] = 14'b00000000111000;
	assign font[15][63] = 14'b00000000111000;
	assign font[16][63] = 14'b00000000111000;
	assign font[17][63] = 14'b00000011100000;
	assign font[18][63] = 14'b00000011100000;
	assign font[19][63] = 14'b00000111000000;
	assign font[20][63] = 14'b00000111000000;
	assign font[21][63] = 14'b00000111000000;
	assign font[22][63] = 14'b00000000000000;
	assign font[23][63] = 14'b00000000000000;
	assign font[24][63] = 14'b00000000000000;
	assign font[25][63] = 14'b00000111000000;
	assign font[26][63] = 14'b00000111000000;
	assign font[27][63] = 14'b00000000000000;
	assign font[28][63] = 14'b00000000000000;
	assign font[29][63] = 14'b00000000000000;
	assign font[30][63] = 14'b00000000000000;
	assign font[31][63] = 14'b00000000000000;

	assign font[0][64] = 14'b00000000000000;
	assign font[1][64] = 14'b00000000000000;
	assign font[2][64] = 14'b00000000000000;
	assign font[3][64] = 14'b00000000000000;
	assign font[4][64] = 14'b00000000000000;
	assign font[5][64] = 14'b00000000000000;
	assign font[6][64] = 14'b00000111111000;
	assign font[7][64] = 14'b00000111111000;
	assign font[8][64] = 14'b00000100011000;
	assign font[9][64] = 14'b00011100011100;
	assign font[10][64] = 14'b00011100011100;
	assign font[11][64] = 14'b00111011111110;
	assign font[12][64] = 14'b00111011111110;
	assign font[13][64] = 14'b00111011111110;
	assign font[14][64] = 14'b00111011001110;
	assign font[15][64] = 14'b00111011001110;
	assign font[16][64] = 14'b00111011001110;
	assign font[17][64] = 14'b00111011001110;
	assign font[18][64] = 14'b00111011001110;
	assign font[19][64] = 14'b00111001111100;
	assign font[20][64] = 14'b00111001111100;
	assign font[21][64] = 14'b00011100000000;
	assign font[22][64] = 14'b00011100000000;
	assign font[23][64] = 14'b00011100000000;
	assign font[24][64] = 14'b00011100000000;
	assign font[25][64] = 14'b00000111111100;
	assign font[26][64] = 14'b00000111111100;
	assign font[27][64] = 14'b00000000000000;
	assign font[28][64] = 14'b00000000000000;
	assign font[29][64] = 14'b00000000000000;
	assign font[30][64] = 14'b00000000000000;
	assign font[31][64] = 14'b00000000000000;

	assign font[0][65] = 14'b00000000000000;
	assign font[1][65] = 14'b00000000000000;
	assign font[2][65] = 14'b00000000000000;
	assign font[3][65] = 14'b00000000000000;
	assign font[4][65] = 14'b00000000000000;
	assign font[5][65] = 14'b00000000000000;
	assign font[6][65] = 14'b00000000000000;
	assign font[7][65] = 14'b00000000000000;
	assign font[8][65] = 14'b00000000000000;
	assign font[9][65] = 14'b00000111100000;
	assign font[10][65] = 14'b00000111100000;
	assign font[11][65] = 14'b00000111110000;
	assign font[12][65] = 14'b00000111110000;
	assign font[13][65] = 14'b00000111110000;
	assign font[14][65] = 14'b00001100111000;
	assign font[15][65] = 14'b00001100111000;
	assign font[16][65] = 14'b00001100111100;
	assign font[17][65] = 14'b00011000011100;
	assign font[18][65] = 14'b00011000011100;
	assign font[19][65] = 14'b00011111111100;
	assign font[20][65] = 14'b00011111111100;
	assign font[21][65] = 14'b00011000001100;
	assign font[22][65] = 14'b00111000001110;
	assign font[23][65] = 14'b00111000001110;
	assign font[24][65] = 14'b00111000001110;
	assign font[25][65] = 14'b00111000001110;
	assign font[26][65] = 14'b00111000001110;
	assign font[27][65] = 14'b00000000000000;
	assign font[28][65] = 14'b00000000000000;
	assign font[29][65] = 14'b00000000000000;
	assign font[30][65] = 14'b00000000000000;
	assign font[31][65] = 14'b00000000000000;

	assign font[0][66] = 14'b00000000000000;
	assign font[1][66] = 14'b00000000000000;
	assign font[2][66] = 14'b00000000000000;
	assign font[3][66] = 14'b00000000000000;
	assign font[4][66] = 14'b00000000000000;
	assign font[5][66] = 14'b00000000000000;
	assign font[6][66] = 14'b00000000000000;
	assign font[7][66] = 14'b00000000000000;
	assign font[8][66] = 14'b00000000000000;
	assign font[9][66] = 14'b00111111111100;
	assign font[10][66] = 14'b00111111111100;
	assign font[11][66] = 14'b00111000001110;
	assign font[12][66] = 14'b00111000001110;
	assign font[13][66] = 14'b00111000001110;
	assign font[14][66] = 14'b00111000001110;
	assign font[15][66] = 14'b00111000001110;
	assign font[16][66] = 14'b00111000001110;
	assign font[17][66] = 14'b00111111111000;
	assign font[18][66] = 14'b00111111111000;
	assign font[19][66] = 14'b00111000001110;
	assign font[20][66] = 14'b00111000001110;
	assign font[21][66] = 14'b00111000001110;
	assign font[22][66] = 14'b00111000001110;
	assign font[23][66] = 14'b00111000001110;
	assign font[24][66] = 14'b00111000001100;
	assign font[25][66] = 14'b00111111111100;
	assign font[26][66] = 14'b00111111111100;
	assign font[27][66] = 14'b00000000000000;
	assign font[28][66] = 14'b00000000000000;
	assign font[29][66] = 14'b00000000000000;
	assign font[30][66] = 14'b00000000000000;
	assign font[31][66] = 14'b00000000000000;

	assign font[0][67] = 14'b00000000000000;
	assign font[1][67] = 14'b00000000000000;
	assign font[2][67] = 14'b00000000000000;
	assign font[3][67] = 14'b00000000000000;
	assign font[4][67] = 14'b00000000000000;
	assign font[5][67] = 14'b00000000000000;
	assign font[6][67] = 14'b00000000000000;
	assign font[7][67] = 14'b00000000000000;
	assign font[8][67] = 14'b00000000000000;
	assign font[9][67] = 14'b00000111111000;
	assign font[10][67] = 14'b00000111111000;
	assign font[11][67] = 14'b00000100001000;
	assign font[12][67] = 14'b00011100001110;
	assign font[13][67] = 14'b00011100001110;
	assign font[14][67] = 14'b00111000000000;
	assign font[15][67] = 14'b00111000000000;
	assign font[16][67] = 14'b00111000000000;
	assign font[17][67] = 14'b00111000000000;
	assign font[18][67] = 14'b00111000000000;
	assign font[19][67] = 14'b00111000000000;
	assign font[20][67] = 14'b00111000000000;
	assign font[21][67] = 14'b00111000000000;
	assign font[22][67] = 14'b00011100001110;
	assign font[23][67] = 14'b00011100001110;
	assign font[24][67] = 14'b00000100001000;
	assign font[25][67] = 14'b00000111111000;
	assign font[26][67] = 14'b00000111111000;
	assign font[27][67] = 14'b00000000000000;
	assign font[28][67] = 14'b00000000000000;
	assign font[29][67] = 14'b00000000000000;
	assign font[30][67] = 14'b00000000000000;
	assign font[31][67] = 14'b00000000000000;

	assign font[0][68] = 14'b00000000000000;
	assign font[1][68] = 14'b00000000000000;
	assign font[2][68] = 14'b00000000000000;
	assign font[3][68] = 14'b00000000000000;
	assign font[4][68] = 14'b00000000000000;
	assign font[5][68] = 14'b00000000000000;
	assign font[6][68] = 14'b00000000000000;
	assign font[7][68] = 14'b00000000000000;
	assign font[8][68] = 14'b00000000000000;
	assign font[9][68] = 14'b00111111110000;
	assign font[10][68] = 14'b00111111110000;
	assign font[11][68] = 14'b00111000011100;
	assign font[12][68] = 14'b00111000011100;
	assign font[13][68] = 14'b00111000011100;
	assign font[14][68] = 14'b00111000001110;
	assign font[15][68] = 14'b00111000001110;
	assign font[16][68] = 14'b00111000001110;
	assign font[17][68] = 14'b00111000001110;
	assign font[18][68] = 14'b00111000001110;
	assign font[19][68] = 14'b00111000001110;
	assign font[20][68] = 14'b00111000001110;
	assign font[21][68] = 14'b00111000001110;
	assign font[22][68] = 14'b00111000011100;
	assign font[23][68] = 14'b00111000011100;
	assign font[24][68] = 14'b00111000010000;
	assign font[25][68] = 14'b00111111110000;
	assign font[26][68] = 14'b00111111110000;
	assign font[27][68] = 14'b00000000000000;
	assign font[28][68] = 14'b00000000000000;
	assign font[29][68] = 14'b00000000000000;
	assign font[30][68] = 14'b00000000000000;
	assign font[31][68] = 14'b00000000000000;

	assign font[0][69] = 14'b00000000000000;
	assign font[1][69] = 14'b00000000000000;
	assign font[2][69] = 14'b00000000000000;
	assign font[3][69] = 14'b00000000000000;
	assign font[4][69] = 14'b00000000000000;
	assign font[5][69] = 14'b00000000000000;
	assign font[6][69] = 14'b00000000000000;
	assign font[7][69] = 14'b00000000000000;
	assign font[8][69] = 14'b00000000000000;
	assign font[9][69] = 14'b00011111111000;
	assign font[10][69] = 14'b00011111111000;
	assign font[11][69] = 14'b00011100000000;
	assign font[12][69] = 14'b00011100000000;
	assign font[13][69] = 14'b00011100000000;
	assign font[14][69] = 14'b00011100000000;
	assign font[15][69] = 14'b00011100000000;
	assign font[16][69] = 14'b00011100000000;
	assign font[17][69] = 14'b00011111111000;
	assign font[18][69] = 14'b00011111111000;
	assign font[19][69] = 14'b00011100000000;
	assign font[20][69] = 14'b00011100000000;
	assign font[21][69] = 14'b00011100000000;
	assign font[22][69] = 14'b00011100000000;
	assign font[23][69] = 14'b00011100000000;
	assign font[24][69] = 14'b00011100000000;
	assign font[25][69] = 14'b00011111111000;
	assign font[26][69] = 14'b00011111111000;
	assign font[27][69] = 14'b00000000000000;
	assign font[28][69] = 14'b00000000000000;
	assign font[29][69] = 14'b00000000000000;
	assign font[30][69] = 14'b00000000000000;
	assign font[31][69] = 14'b00000000000000;

	assign font[0][70] = 14'b00000000000000;
	assign font[1][70] = 14'b00000000000000;
	assign font[2][70] = 14'b00000000000000;
	assign font[3][70] = 14'b00000000000000;
	assign font[4][70] = 14'b00000000000000;
	assign font[5][70] = 14'b00000000000000;
	assign font[6][70] = 14'b00000000000000;
	assign font[7][70] = 14'b00000000000000;
	assign font[8][70] = 14'b00000000000000;
	assign font[9][70] = 14'b00011111111000;
	assign font[10][70] = 14'b00011111111000;
	assign font[11][70] = 14'b00011100000000;
	assign font[12][70] = 14'b00011100000000;
	assign font[13][70] = 14'b00011100000000;
	assign font[14][70] = 14'b00011100000000;
	assign font[15][70] = 14'b00011100000000;
	assign font[16][70] = 14'b00011100000000;
	assign font[17][70] = 14'b00011111111000;
	assign font[18][70] = 14'b00011111111000;
	assign font[19][70] = 14'b00011100000000;
	assign font[20][70] = 14'b00011100000000;
	assign font[21][70] = 14'b00011100000000;
	assign font[22][70] = 14'b00011100000000;
	assign font[23][70] = 14'b00011100000000;
	assign font[24][70] = 14'b00011100000000;
	assign font[25][70] = 14'b00011100000000;
	assign font[26][70] = 14'b00011100000000;
	assign font[27][70] = 14'b00000000000000;
	assign font[28][70] = 14'b00000000000000;
	assign font[29][70] = 14'b00000000000000;
	assign font[30][70] = 14'b00000000000000;
	assign font[31][70] = 14'b00000000000000;

	assign font[0][71] = 14'b00000000000000;
	assign font[1][71] = 14'b00000000000000;
	assign font[2][71] = 14'b00000000000000;
	assign font[3][71] = 14'b00000000000000;
	assign font[4][71] = 14'b00000000000000;
	assign font[5][71] = 14'b00000000000000;
	assign font[6][71] = 14'b00000000000000;
	assign font[7][71] = 14'b00000000000000;
	assign font[8][71] = 14'b00000000000000;
	assign font[9][71] = 14'b00000111111000;
	assign font[10][71] = 14'b00000111111000;
	assign font[11][71] = 14'b00000100001000;
	assign font[12][71] = 14'b00011100001110;
	assign font[13][71] = 14'b00011100001110;
	assign font[14][71] = 14'b00111000000000;
	assign font[15][71] = 14'b00111000000000;
	assign font[16][71] = 14'b00111000000000;
	assign font[17][71] = 14'b00111000111110;
	assign font[18][71] = 14'b00111000111110;
	assign font[19][71] = 14'b00111000111110;
	assign font[20][71] = 14'b00111000001110;
	assign font[21][71] = 14'b00111000001110;
	assign font[22][71] = 14'b00011100001110;
	assign font[23][71] = 14'b00011100001110;
	assign font[24][71] = 14'b00011100001110;
	assign font[25][71] = 14'b00000111111000;
	assign font[26][71] = 14'b00000111111000;
	assign font[27][71] = 14'b00000000000000;
	assign font[28][71] = 14'b00000000000000;
	assign font[29][71] = 14'b00000000000000;
	assign font[30][71] = 14'b00000000000000;
	assign font[31][71] = 14'b00000000000000;

	assign font[0][72] = 14'b00000000000000;
	assign font[1][72] = 14'b00000000000000;
	assign font[2][72] = 14'b00000000000000;
	assign font[3][72] = 14'b00000000000000;
	assign font[4][72] = 14'b00000000000000;
	assign font[5][72] = 14'b00000000000000;
	assign font[6][72] = 14'b00000000000000;
	assign font[7][72] = 14'b00000000000000;
	assign font[8][72] = 14'b00000000000000;
	assign font[9][72] = 14'b00111000001110;
	assign font[10][72] = 14'b00111000001110;
	assign font[11][72] = 14'b00111000001110;
	assign font[12][72] = 14'b00111000001110;
	assign font[13][72] = 14'b00111000001110;
	assign font[14][72] = 14'b00111000001110;
	assign font[15][72] = 14'b00111000001110;
	assign font[16][72] = 14'b00111000001110;
	assign font[17][72] = 14'b00111111111110;
	assign font[18][72] = 14'b00111111111110;
	assign font[19][72] = 14'b00111000001110;
	assign font[20][72] = 14'b00111000001110;
	assign font[21][72] = 14'b00111000001110;
	assign font[22][72] = 14'b00111000001110;
	assign font[23][72] = 14'b00111000001110;
	assign font[24][72] = 14'b00111000001110;
	assign font[25][72] = 14'b00111000001110;
	assign font[26][72] = 14'b00111000001110;
	assign font[27][72] = 14'b00000000000000;
	assign font[28][72] = 14'b00000000000000;
	assign font[29][72] = 14'b00000000000000;
	assign font[30][72] = 14'b00000000000000;
	assign font[31][72] = 14'b00000000000000;

	assign font[0][73] = 14'b00000000000000;
	assign font[1][73] = 14'b00000000000000;
	assign font[2][73] = 14'b00000000000000;
	assign font[3][73] = 14'b00000000000000;
	assign font[4][73] = 14'b00000000000000;
	assign font[5][73] = 14'b00000000000000;
	assign font[6][73] = 14'b00000000000000;
	assign font[7][73] = 14'b00000000000000;
	assign font[8][73] = 14'b00000000000000;
	assign font[9][73] = 14'b00001111110000;
	assign font[10][73] = 14'b00001111110000;
	assign font[11][73] = 14'b00000011100000;
	assign font[12][73] = 14'b00000011100000;
	assign font[13][73] = 14'b00000011100000;
	assign font[14][73] = 14'b00000011100000;
	assign font[15][73] = 14'b00000011100000;
	assign font[16][73] = 14'b00000011100000;
	assign font[17][73] = 14'b00000011100000;
	assign font[18][73] = 14'b00000011100000;
	assign font[19][73] = 14'b00000011100000;
	assign font[20][73] = 14'b00000011100000;
	assign font[21][73] = 14'b00000011100000;
	assign font[22][73] = 14'b00000011100000;
	assign font[23][73] = 14'b00000011100000;
	assign font[24][73] = 14'b00000011100000;
	assign font[25][73] = 14'b00001111110000;
	assign font[26][73] = 14'b00001111110000;
	assign font[27][73] = 14'b00000000000000;
	assign font[28][73] = 14'b00000000000000;
	assign font[29][73] = 14'b00000000000000;
	assign font[30][73] = 14'b00000000000000;
	assign font[31][73] = 14'b00000000000000;

	assign font[0][74] = 14'b00000000000000;
	assign font[1][74] = 14'b00000000000000;
	assign font[2][74] = 14'b00000000000000;
	assign font[3][74] = 14'b00000000000000;
	assign font[4][74] = 14'b00000000000000;
	assign font[5][74] = 14'b00000000000000;
	assign font[6][74] = 14'b00000000000000;
	assign font[7][74] = 14'b00000000000000;
	assign font[8][74] = 14'b00000000000000;
	assign font[9][74] = 14'b00000011111100;
	assign font[10][74] = 14'b00000011111100;
	assign font[11][74] = 14'b00000000111000;
	assign font[12][74] = 14'b00000000111000;
	assign font[13][74] = 14'b00000000111000;
	assign font[14][74] = 14'b00000000111000;
	assign font[15][74] = 14'b00000000111000;
	assign font[16][74] = 14'b00000000111000;
	assign font[17][74] = 14'b00000000111000;
	assign font[18][74] = 14'b00000000111000;
	assign font[19][74] = 14'b00000000111000;
	assign font[20][74] = 14'b00000000111000;
	assign font[21][74] = 14'b00000000111000;
	assign font[22][74] = 14'b00111000111000;
	assign font[23][74] = 14'b00111000111000;
	assign font[24][74] = 14'b00111000111000;
	assign font[25][74] = 14'b00001111110000;
	assign font[26][74] = 14'b00001111110000;
	assign font[27][74] = 14'b00000000000000;
	assign font[28][74] = 14'b00000000000000;
	assign font[29][74] = 14'b00000000000000;
	assign font[30][74] = 14'b00000000000000;
	assign font[31][74] = 14'b00000000000000;

	assign font[0][75] = 14'b00000000000000;
	assign font[1][75] = 14'b00000000000000;
	assign font[2][75] = 14'b00000000000000;
	assign font[3][75] = 14'b00000000000000;
	assign font[4][75] = 14'b00000000000000;
	assign font[5][75] = 14'b00000000000000;
	assign font[6][75] = 14'b00000000000000;
	assign font[7][75] = 14'b00000000000000;
	assign font[8][75] = 14'b00000000000000;
	assign font[9][75] = 14'b00111000011100;
	assign font[10][75] = 14'b00111000011100;
	assign font[11][75] = 14'b00111000011000;
	assign font[12][75] = 14'b00111000111000;
	assign font[13][75] = 14'b00111000111000;
	assign font[14][75] = 14'b00111011100000;
	assign font[15][75] = 14'b00111011100000;
	assign font[16][75] = 14'b00111011000000;
	assign font[17][75] = 14'b00111111000000;
	assign font[18][75] = 14'b00111111000000;
	assign font[19][75] = 14'b00111011100000;
	assign font[20][75] = 14'b00111011100000;
	assign font[21][75] = 14'b00111011100000;
	assign font[22][75] = 14'b00111000111000;
	assign font[23][75] = 14'b00111000111000;
	assign font[24][75] = 14'b00111000011100;
	assign font[25][75] = 14'b00111000011100;
	assign font[26][75] = 14'b00111000011100;
	assign font[27][75] = 14'b00000000000000;
	assign font[28][75] = 14'b00000000000000;
	assign font[29][75] = 14'b00000000000000;
	assign font[30][75] = 14'b00000000000000;
	assign font[31][75] = 14'b00000000000000;

	assign font[0][76] = 14'b00000000000000;
	assign font[1][76] = 14'b00000000000000;
	assign font[2][76] = 14'b00000000000000;
	assign font[3][76] = 14'b00000000000000;
	assign font[4][76] = 14'b00000000000000;
	assign font[5][76] = 14'b00000000000000;
	assign font[6][76] = 14'b00000000000000;
	assign font[7][76] = 14'b00000000000000;
	assign font[8][76] = 14'b00000000000000;
	assign font[9][76] = 14'b00111000000000;
	assign font[10][76] = 14'b00111000000000;
	assign font[11][76] = 14'b00111000000000;
	assign font[12][76] = 14'b00111000000000;
	assign font[13][76] = 14'b00111000000000;
	assign font[14][76] = 14'b00111000000000;
	assign font[15][76] = 14'b00111000000000;
	assign font[16][76] = 14'b00111000000000;
	assign font[17][76] = 14'b00111000000000;
	assign font[18][76] = 14'b00111000000000;
	assign font[19][76] = 14'b00111000000000;
	assign font[20][76] = 14'b00111000000000;
	assign font[21][76] = 14'b00111000000000;
	assign font[22][76] = 14'b00111000000000;
	assign font[23][76] = 14'b00111000000000;
	assign font[24][76] = 14'b00111000000000;
	assign font[25][76] = 14'b00111111111000;
	assign font[26][76] = 14'b00111111111000;
	assign font[27][76] = 14'b00000000000000;
	assign font[28][76] = 14'b00000000000000;
	assign font[29][76] = 14'b00000000000000;
	assign font[30][76] = 14'b00000000000000;
	assign font[31][76] = 14'b00000000000000;

	assign font[0][77] = 14'b00000000000000;
	assign font[1][77] = 14'b00000000000000;
	assign font[2][77] = 14'b00000000000000;
	assign font[3][77] = 14'b00000000000000;
	assign font[4][77] = 14'b00000000000000;
	assign font[5][77] = 14'b00000000000000;
	assign font[6][77] = 14'b00000000000000;
	assign font[7][77] = 14'b00000000000000;
	assign font[8][77] = 14'b00000000000000;
	assign font[9][77] = 14'b00111100011110;
	assign font[10][77] = 14'b00111100011110;
	assign font[11][77] = 14'b00111110111110;
	assign font[12][77] = 14'b00111110111110;
	assign font[13][77] = 14'b00111110111110;
	assign font[14][77] = 14'b00111010101110;
	assign font[15][77] = 14'b00111010101110;
	assign font[16][77] = 14'b00111011101110;
	assign font[17][77] = 14'b00111011101110;
	assign font[18][77] = 14'b00111011101110;
	assign font[19][77] = 14'b00111011001110;
	assign font[20][77] = 14'b00111011001110;
	assign font[21][77] = 14'b00111001001110;
	assign font[22][77] = 14'b00111011001110;
	assign font[23][77] = 14'b00111011001110;
	assign font[24][77] = 14'b00111000001110;
	assign font[25][77] = 14'b00111000001110;
	assign font[26][77] = 14'b00111000001110;
	assign font[27][77] = 14'b00000000000000;
	assign font[28][77] = 14'b00000000000000;
	assign font[29][77] = 14'b00000000000000;
	assign font[30][77] = 14'b00000000000000;
	assign font[31][77] = 14'b00000000000000;

	assign font[0][78] = 14'b00000000000000;
	assign font[1][78] = 14'b00000000000000;
	assign font[2][78] = 14'b00000000000000;
	assign font[3][78] = 14'b00000000000000;
	assign font[4][78] = 14'b00000000000000;
	assign font[5][78] = 14'b00000000000000;
	assign font[6][78] = 14'b00000000000000;
	assign font[7][78] = 14'b00000000000000;
	assign font[8][78] = 14'b00000000000000;
	assign font[9][78] = 14'b00111000001110;
	assign font[10][78] = 14'b00111000001110;
	assign font[11][78] = 14'b00111100001110;
	assign font[12][78] = 14'b00111100001110;
	assign font[13][78] = 14'b00111100001110;
	assign font[14][78] = 14'b00111111001110;
	assign font[15][78] = 14'b00111111001110;
	assign font[16][78] = 14'b00111111001110;
	assign font[17][78] = 14'b00111011101110;
	assign font[18][78] = 14'b00111011101110;
	assign font[19][78] = 14'b00111001111110;
	assign font[20][78] = 14'b00111001111110;
	assign font[21][78] = 14'b00111001111110;
	assign font[22][78] = 14'b00111000111110;
	assign font[23][78] = 14'b00111000111110;
	assign font[24][78] = 14'b00111000001110;
	assign font[25][78] = 14'b00111000001110;
	assign font[26][78] = 14'b00111000001110;
	assign font[27][78] = 14'b00000000000000;
	assign font[28][78] = 14'b00000000000000;
	assign font[29][78] = 14'b00000000000000;
	assign font[30][78] = 14'b00000000000000;
	assign font[31][78] = 14'b00000000000000;

	assign font[0][79] = 14'b00000000000000;
	assign font[1][79] = 14'b00000000000000;
	assign font[2][79] = 14'b00000000000000;
	assign font[3][79] = 14'b00000000000000;
	assign font[4][79] = 14'b00000000000000;
	assign font[5][79] = 14'b00000000000000;
	assign font[6][79] = 14'b00000000000000;
	assign font[7][79] = 14'b00000000000000;
	assign font[8][79] = 14'b00000000000000;
	assign font[9][79] = 14'b00001111110000;
	assign font[10][79] = 14'b00001111110000;
	assign font[11][79] = 14'b00011100011100;
	assign font[12][79] = 14'b00011100011100;
	assign font[13][79] = 14'b00011100011100;
	assign font[14][79] = 14'b00111000001110;
	assign font[15][79] = 14'b00111000001110;
	assign font[16][79] = 14'b00111000001110;
	assign font[17][79] = 14'b00111000001110;
	assign font[18][79] = 14'b00111000001110;
	assign font[19][79] = 14'b00111000001110;
	assign font[20][79] = 14'b00111000001110;
	assign font[21][79] = 14'b00111000001110;
	assign font[22][79] = 14'b00011100011100;
	assign font[23][79] = 14'b00011100011100;
	assign font[24][79] = 14'b00001100010000;
	assign font[25][79] = 14'b00001111110000;
	assign font[26][79] = 14'b00001111110000;
	assign font[27][79] = 14'b00000000000000;
	assign font[28][79] = 14'b00000000000000;
	assign font[29][79] = 14'b00000000000000;
	assign font[30][79] = 14'b00000000000000;
	assign font[31][79] = 14'b00000000000000;

	assign font[0][80] = 14'b00000000000000;
	assign font[1][80] = 14'b00000000000000;
	assign font[2][80] = 14'b00000000000000;
	assign font[3][80] = 14'b00000000000000;
	assign font[4][80] = 14'b00000000000000;
	assign font[5][80] = 14'b00000000000000;
	assign font[6][80] = 14'b00000000000000;
	assign font[7][80] = 14'b00000000000000;
	assign font[8][80] = 14'b00000000000000;
	assign font[9][80] = 14'b00111111110000;
	assign font[10][80] = 14'b00111111110000;
	assign font[11][80] = 14'b00111000011100;
	assign font[12][80] = 14'b00111000011100;
	assign font[13][80] = 14'b00111000011100;
	assign font[14][80] = 14'b00111000011100;
	assign font[15][80] = 14'b00111000011100;
	assign font[16][80] = 14'b00111000010000;
	assign font[17][80] = 14'b00111111110000;
	assign font[18][80] = 14'b00111111110000;
	assign font[19][80] = 14'b00111000000000;
	assign font[20][80] = 14'b00111000000000;
	assign font[21][80] = 14'b00111000000000;
	assign font[22][80] = 14'b00111000000000;
	assign font[23][80] = 14'b00111000000000;
	assign font[24][80] = 14'b00111000000000;
	assign font[25][80] = 14'b00111000000000;
	assign font[26][80] = 14'b00111000000000;
	assign font[27][80] = 14'b00000000000000;
	assign font[28][80] = 14'b00000000000000;
	assign font[29][80] = 14'b00000000000000;
	assign font[30][80] = 14'b00000000000000;
	assign font[31][80] = 14'b00000000000000;

	assign font[0][81] = 14'b00000000000000;
	assign font[1][81] = 14'b00000000000000;
	assign font[2][81] = 14'b00000000000000;
	assign font[3][81] = 14'b00000000000000;
	assign font[4][81] = 14'b00000000000000;
	assign font[5][81] = 14'b00000000000000;
	assign font[6][81] = 14'b00000000000000;
	assign font[7][81] = 14'b00000000000000;
	assign font[8][81] = 14'b00000000000000;
	assign font[9][81] = 14'b00001111110000;
	assign font[10][81] = 14'b00001111110000;
	assign font[11][81] = 14'b00011100011100;
	assign font[12][81] = 14'b00011100011100;
	assign font[13][81] = 14'b00011100011100;
	assign font[14][81] = 14'b00111000001110;
	assign font[15][81] = 14'b00111000001110;
	assign font[16][81] = 14'b00111000001110;
	assign font[17][81] = 14'b00111000001110;
	assign font[18][81] = 14'b00111000001110;
	assign font[19][81] = 14'b00111011101110;
	assign font[20][81] = 14'b00111011101110;
	assign font[21][81] = 14'b00111011101110;
	assign font[22][81] = 14'b00011101111100;
	assign font[23][81] = 14'b00011101111100;
	assign font[24][81] = 14'b00001101110000;
	assign font[25][81] = 14'b00001111110000;
	assign font[26][81] = 14'b00001111110000;
	assign font[27][81] = 14'b00000000011000;
	assign font[28][81] = 14'b00000000011000;
	assign font[29][81] = 14'b00000000001100;
	assign font[30][81] = 14'b00000000001100;
	assign font[31][81] = 14'b00000000001100;

	assign font[0][82] = 14'b00000000000000;
	assign font[1][82] = 14'b00000000000000;
	assign font[2][82] = 14'b00000000000000;
	assign font[3][82] = 14'b00000000000000;
	assign font[4][82] = 14'b00000000000000;
	assign font[5][82] = 14'b00000000000000;
	assign font[6][82] = 14'b00000000000000;
	assign font[7][82] = 14'b00000000000000;
	assign font[8][82] = 14'b00000000000000;
	assign font[9][82] = 14'b00111111111000;
	assign font[10][82] = 14'b00111111111000;
	assign font[11][82] = 14'b00111000011000;
	assign font[12][82] = 14'b00111000011110;
	assign font[13][82] = 14'b00111000011110;
	assign font[14][82] = 14'b00111000011100;
	assign font[15][82] = 14'b00111000011100;
	assign font[16][82] = 14'b00111000011100;
	assign font[17][82] = 14'b00111111110000;
	assign font[18][82] = 14'b00111111110000;
	assign font[19][82] = 14'b00111000111000;
	assign font[20][82] = 14'b00111000111000;
	assign font[21][82] = 14'b00111000111000;
	assign font[22][82] = 14'b00111000011100;
	assign font[23][82] = 14'b00111000011100;
	assign font[24][82] = 14'b00111000011100;
	assign font[25][82] = 14'b00111000001110;
	assign font[26][82] = 14'b00111000001110;
	assign font[27][82] = 14'b00000000000000;
	assign font[28][82] = 14'b00000000000000;
	assign font[29][82] = 14'b00000000000000;
	assign font[30][82] = 14'b00000000000000;
	assign font[31][82] = 14'b00000000000000;

	assign font[0][83] = 14'b00000000000000;
	assign font[1][83] = 14'b00000000000000;
	assign font[2][83] = 14'b00000000000000;
	assign font[3][83] = 14'b00000000000000;
	assign font[4][83] = 14'b00000000000000;
	assign font[5][83] = 14'b00000000000000;
	assign font[6][83] = 14'b00000000000000;
	assign font[7][83] = 14'b00000000000000;
	assign font[8][83] = 14'b00000000000000;
	assign font[9][83] = 14'b00001111111000;
	assign font[10][83] = 14'b00001111111000;
	assign font[11][83] = 14'b00001000001000;
	assign font[12][83] = 14'b00111000001110;
	assign font[13][83] = 14'b00111000001110;
	assign font[14][83] = 14'b00111000000000;
	assign font[15][83] = 14'b00111000000000;
	assign font[16][83] = 14'b00111000000000;
	assign font[17][83] = 14'b00001111111000;
	assign font[18][83] = 14'b00001111111000;
	assign font[19][83] = 14'b00000000001110;
	assign font[20][83] = 14'b00000000001110;
	assign font[21][83] = 14'b00000000001110;
	assign font[22][83] = 14'b00111000001110;
	assign font[23][83] = 14'b00111000001110;
	assign font[24][83] = 14'b00001000001000;
	assign font[25][83] = 14'b00001111111000;
	assign font[26][83] = 14'b00001111111000;
	assign font[27][83] = 14'b00000000000000;
	assign font[28][83] = 14'b00000000000000;
	assign font[29][83] = 14'b00000000000000;
	assign font[30][83] = 14'b00000000000000;
	assign font[31][83] = 14'b00000000000000;

	assign font[0][84] = 14'b00000000000000;
	assign font[1][84] = 14'b00000000000000;
	assign font[2][84] = 14'b00000000000000;
	assign font[3][84] = 14'b00000000000000;
	assign font[4][84] = 14'b00000000000000;
	assign font[5][84] = 14'b00000000000000;
	assign font[6][84] = 14'b00000000000000;
	assign font[7][84] = 14'b00000000000000;
	assign font[8][84] = 14'b00000000000000;
	assign font[9][84] = 14'b00111111111100;
	assign font[10][84] = 14'b00011111111100;
	assign font[11][84] = 14'b00000011100000;
	assign font[12][84] = 14'b00000011100000;
	assign font[13][84] = 14'b00000011100000;
	assign font[14][84] = 14'b00000011100000;
	assign font[15][84] = 14'b00000011100000;
	assign font[16][84] = 14'b00000011100000;
	assign font[17][84] = 14'b00000011100000;
	assign font[18][84] = 14'b00000011100000;
	assign font[19][84] = 14'b00000011100000;
	assign font[20][84] = 14'b00000011100000;
	assign font[21][84] = 14'b00000011100000;
	assign font[22][84] = 14'b00000011100000;
	assign font[23][84] = 14'b00000011100000;
	assign font[24][84] = 14'b00000011100000;
	assign font[25][84] = 14'b00000011100000;
	assign font[26][84] = 14'b00000011100000;
	assign font[27][84] = 14'b00000000000000;
	assign font[28][84] = 14'b00000000000000;
	assign font[29][84] = 14'b00000000000000;
	assign font[30][84] = 14'b00000000000000;
	assign font[31][84] = 14'b00000000000000;

	assign font[0][85] = 14'b00000000000000;
	assign font[1][85] = 14'b00000000000000;
	assign font[2][85] = 14'b00000000000000;
	assign font[3][85] = 14'b00000000000000;
	assign font[4][85] = 14'b00000000000000;
	assign font[5][85] = 14'b00000000000000;
	assign font[6][85] = 14'b00000000000000;
	assign font[7][85] = 14'b00000000000000;
	assign font[8][85] = 14'b00000000000000;
	assign font[9][85] = 14'b00111000001110;
	assign font[10][85] = 14'b00111000001110;
	assign font[11][85] = 14'b00111000001110;
	assign font[12][85] = 14'b00111000001110;
	assign font[13][85] = 14'b00111000001110;
	assign font[14][85] = 14'b00111000001110;
	assign font[15][85] = 14'b00111000001110;
	assign font[16][85] = 14'b00111000001110;
	assign font[17][85] = 14'b00111000001110;
	assign font[18][85] = 14'b00111000001110;
	assign font[19][85] = 14'b00111000001110;
	assign font[20][85] = 14'b00111000001110;
	assign font[21][85] = 14'b00111000001110;
	assign font[22][85] = 14'b00111000001110;
	assign font[23][85] = 14'b00111000001110;
	assign font[24][85] = 14'b00001000001000;
	assign font[25][85] = 14'b00001111111000;
	assign font[26][85] = 14'b00001111111000;
	assign font[27][85] = 14'b00000000000000;
	assign font[28][85] = 14'b00000000000000;
	assign font[29][85] = 14'b00000000000000;
	assign font[30][85] = 14'b00000000000000;
	assign font[31][85] = 14'b00000000000000;

	assign font[0][86] = 14'b00000000000000;
	assign font[1][86] = 14'b00000000000000;
	assign font[2][86] = 14'b00000000000000;
	assign font[3][86] = 14'b00000000000000;
	assign font[4][86] = 14'b00000000000000;
	assign font[5][86] = 14'b00000000000000;
	assign font[6][86] = 14'b00000000000000;
	assign font[7][86] = 14'b00000000000000;
	assign font[8][86] = 14'b00000000000000;
	assign font[9][86] = 14'b00111000011100;
	assign font[10][86] = 14'b00111000011100;
	assign font[11][86] = 14'b00111000011100;
	assign font[12][86] = 14'b00111000011100;
	assign font[13][86] = 14'b00111000011100;
	assign font[14][86] = 14'b00111000011100;
	assign font[15][86] = 14'b00111000011100;
	assign font[16][86] = 14'b00111000011100;
	assign font[17][86] = 14'b00011100011000;
	assign font[18][86] = 14'b00011100011000;
	assign font[19][86] = 14'b00011110111000;
	assign font[20][86] = 14'b00001110111000;
	assign font[21][86] = 14'b00001110111000;
	assign font[22][86] = 14'b00000111110000;
	assign font[23][86] = 14'b00000111110000;
	assign font[24][86] = 14'b00000111110000;
	assign font[25][86] = 14'b00000011100000;
	assign font[26][86] = 14'b00000011100000;
	assign font[27][86] = 14'b00000000000000;
	assign font[28][86] = 14'b00000000000000;
	assign font[29][86] = 14'b00000000000000;
	assign font[30][86] = 14'b00000000000000;
	assign font[31][86] = 14'b00000000000000;

	assign font[0][87] = 14'b00000000000000;
	assign font[1][87] = 14'b00000000000000;
	assign font[2][87] = 14'b00000000000000;
	assign font[3][87] = 14'b00000000000000;
	assign font[4][87] = 14'b00000000000000;
	assign font[5][87] = 14'b00000000000000;
	assign font[6][87] = 14'b00000000000000;
	assign font[7][87] = 14'b00000000000000;
	assign font[8][87] = 14'b00000000000000;
	assign font[9][87] = 14'b00111011001110;
	assign font[10][87] = 14'b00111011001110;
	assign font[11][87] = 14'b00111011001110;
	assign font[12][87] = 14'b00111011001110;
	assign font[13][87] = 14'b00111011001110;
	assign font[14][87] = 14'b00111011001110;
	assign font[15][87] = 14'b00111011001110;
	assign font[16][87] = 14'b00111011001110;
	assign font[17][87] = 14'b00111011001110;
	assign font[18][87] = 14'b00111011001110;
	assign font[19][87] = 14'b00011011101100;
	assign font[20][87] = 14'b00011011101100;
	assign font[21][87] = 14'b00011011101100;
	assign font[22][87] = 14'b00011110111100;
	assign font[23][87] = 14'b00011110111100;
	assign font[24][87] = 14'b00001100011000;
	assign font[25][87] = 14'b00001100011000;
	assign font[26][87] = 14'b00001100011000;
	assign font[27][87] = 14'b00000000000000;
	assign font[28][87] = 14'b00000000000000;
	assign font[29][87] = 14'b00000000000000;
	assign font[30][87] = 14'b00000000000000;
	assign font[31][87] = 14'b00000000000000;

	assign font[0][88] = 14'b00000000000000;
	assign font[1][88] = 14'b00000000000000;
	assign font[2][88] = 14'b00000000000000;
	assign font[3][88] = 14'b00000000000000;
	assign font[4][88] = 14'b00000000000000;
	assign font[5][88] = 14'b00000000000000;
	assign font[6][88] = 14'b00000000000000;
	assign font[7][88] = 14'b00000000000000;
	assign font[8][88] = 14'b00000000000000;
	assign font[9][88] = 14'b00111000001110;
	assign font[10][88] = 14'b00111000001110;
	assign font[11][88] = 14'b00011100011100;
	assign font[12][88] = 14'b00011100011100;
	assign font[13][88] = 14'b00011100011100;
	assign font[14][88] = 14'b00000110110000;
	assign font[15][88] = 14'b00000110110000;
	assign font[16][88] = 14'b00000110110000;
	assign font[17][88] = 14'b00000111100000;
	assign font[18][88] = 14'b00000111100000;
	assign font[19][88] = 14'b00000110110000;
	assign font[20][88] = 14'b00000110110000;
	assign font[21][88] = 14'b00000110110000;
	assign font[22][88] = 14'b00011100011100;
	assign font[23][88] = 14'b00011100011100;
	assign font[24][88] = 14'b00011000001110;
	assign font[25][88] = 14'b00111000001110;
	assign font[26][88] = 14'b00111000001110;
	assign font[27][88] = 14'b00000000000000;
	assign font[28][88] = 14'b00000000000000;
	assign font[29][88] = 14'b00000000000000;
	assign font[30][88] = 14'b00000000000000;
	assign font[31][88] = 14'b00000000000000;

	assign font[0][89] = 14'b00000000000000;
	assign font[1][89] = 14'b00000000000000;
	assign font[2][89] = 14'b00000000000000;
	assign font[3][89] = 14'b00000000000000;
	assign font[4][89] = 14'b00000000000000;
	assign font[5][89] = 14'b00000000000000;
	assign font[6][89] = 14'b00000000000000;
	assign font[7][89] = 14'b00000000000000;
	assign font[8][89] = 14'b00000000000000;
	assign font[9][89] = 14'b00111000011100;
	assign font[10][89] = 14'b00111000011100;
	assign font[11][89] = 14'b00111000011100;
	assign font[12][89] = 14'b00111000011100;
	assign font[13][89] = 14'b00111000011100;
	assign font[14][89] = 14'b00011100011000;
	assign font[15][89] = 14'b00011100011000;
	assign font[16][89] = 14'b00011100011000;
	assign font[17][89] = 14'b00001111110000;
	assign font[18][89] = 14'b00001111110000;
	assign font[19][89] = 14'b00000011100000;
	assign font[20][89] = 14'b00000011100000;
	assign font[21][89] = 14'b00000011100000;
	assign font[22][89] = 14'b00000011100000;
	assign font[23][89] = 14'b00000011100000;
	assign font[24][89] = 14'b00000011100000;
	assign font[25][89] = 14'b00000011100000;
	assign font[26][89] = 14'b00000011100000;
	assign font[27][89] = 14'b00000000000000;
	assign font[28][89] = 14'b00000000000000;
	assign font[29][89] = 14'b00000000000000;
	assign font[30][89] = 14'b00000000000000;
	assign font[31][89] = 14'b00000000000000;

	assign font[0][90] = 14'b00000000000000;
	assign font[1][90] = 14'b00000000000000;
	assign font[2][90] = 14'b00000000000000;
	assign font[3][90] = 14'b00000000000000;
	assign font[4][90] = 14'b00000000000000;
	assign font[5][90] = 14'b00000000000000;
	assign font[6][90] = 14'b00000000000000;
	assign font[7][90] = 14'b00000000000000;
	assign font[8][90] = 14'b00000000000000;
	assign font[9][90] = 14'b00111111111000;
	assign font[10][90] = 14'b00111111111000;
	assign font[11][90] = 14'b00000000111000;
	assign font[12][90] = 14'b00000000111000;
	assign font[13][90] = 14'b00000000111000;
	assign font[14][90] = 14'b00000001110000;
	assign font[15][90] = 14'b00000001110000;
	assign font[16][90] = 14'b00000001110000;
	assign font[17][90] = 14'b00000011100000;
	assign font[18][90] = 14'b00000011100000;
	assign font[19][90] = 14'b00000011100000;
	assign font[20][90] = 14'b00001110000000;
	assign font[21][90] = 14'b00001110000000;
	assign font[22][90] = 14'b00111000000000;
	assign font[23][90] = 14'b00111000000000;
	assign font[24][90] = 14'b00111000000000;
	assign font[25][90] = 14'b00111111111000;
	assign font[26][90] = 14'b00111111111000;
	assign font[27][90] = 14'b00000000000000;
	assign font[28][90] = 14'b00000000000000;
	assign font[29][90] = 14'b00000000000000;
	assign font[30][90] = 14'b00000000000000;
	assign font[31][90] = 14'b00000000000000;

	assign font[0][91] = 14'b00000000000000;
	assign font[1][91] = 14'b00000000000000;
	assign font[2][91] = 14'b00000000000000;
	assign font[3][91] = 14'b00000000000000;
	assign font[4][91] = 14'b00000000000000;
	assign font[5][91] = 14'b00000000000000;
	assign font[6][91] = 14'b00000000000000;
	assign font[7][91] = 14'b00000111110000;
	assign font[8][91] = 14'b00000111110000;
	assign font[9][91] = 14'b00000111000000;
	assign font[10][91] = 14'b00000111000000;
	assign font[11][91] = 14'b00000111000000;
	assign font[12][91] = 14'b00000111000000;
	assign font[13][91] = 14'b00000111000000;
	assign font[14][91] = 14'b00000111000000;
	assign font[15][91] = 14'b00000111000000;
	assign font[16][91] = 14'b00000111000000;
	assign font[17][91] = 14'b00000111000000;
	assign font[18][91] = 14'b00000111000000;
	assign font[19][91] = 14'b00000111000000;
	assign font[20][91] = 14'b00000111000000;
	assign font[21][91] = 14'b00000111000000;
	assign font[22][91] = 14'b00000111000000;
	assign font[23][91] = 14'b00000111000000;
	assign font[24][91] = 14'b00000111000000;
	assign font[25][91] = 14'b00000111000000;
	assign font[26][91] = 14'b00000111000000;
	assign font[27][91] = 14'b00000111000000;
	assign font[28][91] = 14'b00000111110000;
	assign font[29][91] = 14'b00000111110000;
	assign font[30][91] = 14'b00000000000000;
	assign font[31][91] = 14'b00000000000000;

	assign font[0][92] = 14'b00000000000000;
	assign font[1][92] = 14'b00000000000000;
	assign font[2][92] = 14'b00000000000000;
	assign font[3][92] = 14'b00000000000000;
	assign font[4][92] = 14'b00000000000000;
	assign font[5][92] = 14'b00000000000000;
	assign font[6][92] = 14'b00111000000000;
	assign font[7][92] = 14'b00111000000000;
	assign font[8][92] = 14'b00111000000000;
	assign font[9][92] = 14'b00011100000000;
	assign font[10][92] = 14'b00011100000000;
	assign font[11][92] = 14'b00011100000000;
	assign font[12][92] = 14'b00001110000000;
	assign font[13][92] = 14'b00001110000000;
	assign font[14][92] = 14'b00000111000000;
	assign font[15][92] = 14'b00000111000000;
	assign font[16][92] = 14'b00000111000000;
	assign font[17][92] = 14'b00000011100000;
	assign font[18][92] = 14'b00000011100000;
	assign font[19][92] = 14'b00000011100000;
	assign font[20][92] = 14'b00000011100000;
	assign font[21][92] = 14'b00000011100000;
	assign font[22][92] = 14'b00000000110000;
	assign font[23][92] = 14'b00000000110000;
	assign font[24][92] = 14'b00000000011000;
	assign font[25][92] = 14'b00000000011000;
	assign font[26][92] = 14'b00000000011000;
	assign font[27][92] = 14'b00000000011100;
	assign font[28][92] = 14'b00000000011100;
	assign font[29][92] = 14'b00000000000000;
	assign font[30][92] = 14'b00000000000000;
	assign font[31][92] = 14'b00000000000000;

	assign font[0][93] = 14'b00000000000000;
	assign font[1][93] = 14'b00000000000000;
	assign font[2][93] = 14'b00000000000000;
	assign font[3][93] = 14'b00000000000000;
	assign font[4][93] = 14'b00000000000000;
	assign font[5][93] = 14'b00000000000000;
	assign font[6][93] = 14'b00000000000000;
	assign font[7][93] = 14'b00000111110000;
	assign font[8][93] = 14'b00000111110000;
	assign font[9][93] = 14'b00000001110000;
	assign font[10][93] = 14'b00000001110000;
	assign font[11][93] = 14'b00000001110000;
	assign font[12][93] = 14'b00000001110000;
	assign font[13][93] = 14'b00000001110000;
	assign font[14][93] = 14'b00000001110000;
	assign font[15][93] = 14'b00000001110000;
	assign font[16][93] = 14'b00000001110000;
	assign font[17][93] = 14'b00000001110000;
	assign font[18][93] = 14'b00000001110000;
	assign font[19][93] = 14'b00000001110000;
	assign font[20][93] = 14'b00000001110000;
	assign font[21][93] = 14'b00000001110000;
	assign font[22][93] = 14'b00000001110000;
	assign font[23][93] = 14'b00000001110000;
	assign font[24][93] = 14'b00000001110000;
	assign font[25][93] = 14'b00000001110000;
	assign font[26][93] = 14'b00000001110000;
	assign font[27][93] = 14'b00000001110000;
	assign font[28][93] = 14'b00000111110000;
	assign font[29][93] = 14'b00000111110000;
	assign font[30][93] = 14'b00000000000000;
	assign font[31][93] = 14'b00000000000000;

	assign font[0][94] = 14'b00000000000000;
	assign font[1][94] = 14'b00000000000000;
	assign font[2][94] = 14'b00000000000000;
	assign font[3][94] = 14'b00000000000000;
	assign font[4][94] = 14'b00000000000000;
	assign font[5][94] = 14'b00000000000000;
	assign font[6][94] = 14'b00000000000000;
	assign font[7][94] = 14'b00000000000000;
	assign font[8][94] = 14'b00000000000000;
	assign font[9][94] = 14'b00000111110000;
	assign font[10][94] = 14'b00000111110000;
	assign font[11][94] = 14'b00000111111000;
	assign font[12][94] = 14'b00001110111000;
	assign font[13][94] = 14'b00001110111000;
	assign font[14][94] = 14'b00011100011100;
	assign font[15][94] = 14'b00011100011100;
	assign font[16][94] = 14'b00011100011100;
	assign font[17][94] = 14'b00000000000000;
	assign font[18][94] = 14'b00000000000000;
	assign font[19][94] = 14'b00000000000000;
	assign font[20][94] = 14'b00000000000000;
	assign font[21][94] = 14'b00000000000000;
	assign font[22][94] = 14'b00000000000000;
	assign font[23][94] = 14'b00000000000000;
	assign font[24][94] = 14'b00000000000000;
	assign font[25][94] = 14'b00000000000000;
	assign font[26][94] = 14'b00000000000000;
	assign font[27][94] = 14'b00000000000000;
	assign font[28][94] = 14'b00000000000000;
	assign font[29][94] = 14'b00000000000000;
	assign font[30][94] = 14'b00000000000000;
	assign font[31][94] = 14'b00000000000000;

	assign font[0][95] = 14'b00000000000000;
	assign font[1][95] = 14'b00000000000000;
	assign font[2][95] = 14'b00000000000000;
	assign font[3][95] = 14'b00000000000000;
	assign font[4][95] = 14'b00000000000000;
	assign font[5][95] = 14'b00000000000000;
	assign font[6][95] = 14'b00000000000000;
	assign font[7][95] = 14'b00000000000000;
	assign font[8][95] = 14'b00000000000000;
	assign font[9][95] = 14'b00000000000000;
	assign font[10][95] = 14'b00000000000000;
	assign font[11][95] = 14'b00000000000000;
	assign font[12][95] = 14'b00000000000000;
	assign font[13][95] = 14'b00000000000000;
	assign font[14][95] = 14'b00000000000000;
	assign font[15][95] = 14'b00000000000000;
	assign font[16][95] = 14'b00000000000000;
	assign font[17][95] = 14'b00000000000000;
	assign font[18][95] = 14'b00000000000000;
	assign font[19][95] = 14'b00000000000000;
	assign font[20][95] = 14'b00000000000000;
	assign font[21][95] = 14'b00000000000000;
	assign font[22][95] = 14'b00000000000000;
	assign font[23][95] = 14'b00000000000000;
	assign font[24][95] = 14'b00000000000000;
	assign font[25][95] = 14'b00111111111110;
	assign font[26][95] = 14'b00111111111110;
	assign font[27][95] = 14'b00000000000000;
	assign font[28][95] = 14'b00000000000000;
	assign font[29][95] = 14'b00000000000000;
	assign font[30][95] = 14'b00000000000000;
	assign font[31][95] = 14'b00000000000000;

	assign font[0][96] = 14'b00000000000000;
	assign font[1][96] = 14'b00000000000000;
	assign font[2][96] = 14'b00000000000000;
	assign font[3][96] = 14'b00000000000000;
	assign font[4][96] = 14'b00000000000000;
	assign font[5][96] = 14'b00000000000000;
	assign font[6][96] = 14'b00001110000000;
	assign font[7][96] = 14'b00001110000000;
	assign font[8][96] = 14'b00000010000000;
	assign font[9][96] = 14'b00000011100000;
	assign font[10][96] = 14'b00000011100000;
	assign font[11][96] = 14'b00000000000000;
	assign font[12][96] = 14'b00000000000000;
	assign font[13][96] = 14'b00000000000000;
	assign font[14][96] = 14'b00000000000000;
	assign font[15][96] = 14'b00000000000000;
	assign font[16][96] = 14'b00000000000000;
	assign font[17][96] = 14'b00000000000000;
	assign font[18][96] = 14'b00000000000000;
	assign font[19][96] = 14'b00000000000000;
	assign font[20][96] = 14'b00000000000000;
	assign font[21][96] = 14'b00000000000000;
	assign font[22][96] = 14'b00000000000000;
	assign font[23][96] = 14'b00000000000000;
	assign font[24][96] = 14'b00000000000000;
	assign font[25][96] = 14'b00000000000000;
	assign font[26][96] = 14'b00000000000000;
	assign font[27][96] = 14'b00000000000000;
	assign font[28][96] = 14'b00000000000000;
	assign font[29][96] = 14'b00000000000000;
	assign font[30][96] = 14'b00000000000000;
	assign font[31][96] = 14'b00000000000000;

	assign font[0][97] = 14'b00000000000000;
	assign font[1][97] = 14'b00000000000000;
	assign font[2][97] = 14'b00000000000000;
	assign font[3][97] = 14'b00000000000000;
	assign font[4][97] = 14'b00000000000000;
	assign font[5][97] = 14'b00000000000000;
	assign font[6][97] = 14'b00000000000000;
	assign font[7][97] = 14'b00000000000000;
	assign font[8][97] = 14'b00000000000000;
	assign font[9][97] = 14'b00000000000000;
	assign font[10][97] = 14'b00000000000000;
	assign font[11][97] = 14'b00000000000000;
	assign font[12][97] = 14'b00000000000000;
	assign font[13][97] = 14'b00000000000000;
	assign font[14][97] = 14'b00000111111000;
	assign font[15][97] = 14'b00000111111000;
	assign font[16][97] = 14'b00000000011000;
	assign font[17][97] = 14'b00000000011100;
	assign font[18][97] = 14'b00000000011100;
	assign font[19][97] = 14'b00001111111100;
	assign font[20][97] = 14'b00001111111100;
	assign font[21][97] = 14'b00001111111100;
	assign font[22][97] = 14'b00011100011100;
	assign font[23][97] = 14'b00011100011100;
	assign font[24][97] = 14'b00001111111110;
	assign font[25][97] = 14'b00001111111110;
	assign font[26][97] = 14'b00001111111110;
	assign font[27][97] = 14'b00000000000000;
	assign font[28][97] = 14'b00000000000000;
	assign font[29][97] = 14'b00000000000000;
	assign font[30][97] = 14'b00000000000000;
	assign font[31][97] = 14'b00000000000000;

	assign font[0][98] = 14'b00000000000000;
	assign font[1][98] = 14'b00000000000000;
	assign font[2][98] = 14'b00000000000000;
	assign font[3][98] = 14'b00000000000000;
	assign font[4][98] = 14'b00000000000000;
	assign font[5][98] = 14'b00000000000000;
	assign font[6][98] = 14'b00000000000000;
	assign font[7][98] = 14'b00000000000000;
	assign font[8][98] = 14'b00000000000000;
	assign font[9][98] = 14'b00111000000000;
	assign font[10][98] = 14'b00111000000000;
	assign font[11][98] = 14'b00111000000000;
	assign font[12][98] = 14'b00111000000000;
	assign font[13][98] = 14'b00111000000000;
	assign font[14][98] = 14'b00111111110000;
	assign font[15][98] = 14'b00111111110000;
	assign font[16][98] = 14'b00111100001100;
	assign font[17][98] = 14'b00111100001100;
	assign font[18][98] = 14'b00111100001100;
	assign font[19][98] = 14'b00111000001110;
	assign font[20][98] = 14'b00111000001110;
	assign font[21][98] = 14'b00111000001100;
	assign font[22][98] = 14'b00111000001100;
	assign font[23][98] = 14'b00111000001100;
	assign font[24][98] = 14'b00110000000000;
	assign font[25][98] = 14'b00110111110000;
	assign font[26][98] = 14'b00110111110000;
	assign font[27][98] = 14'b00000000000000;
	assign font[28][98] = 14'b00000000000000;
	assign font[29][98] = 14'b00000000000000;
	assign font[30][98] = 14'b00000000000000;
	assign font[31][98] = 14'b00000000000000;

	assign font[0][99] = 14'b00000000000000;
	assign font[1][99] = 14'b00000000000000;
	assign font[2][99] = 14'b00000000000000;
	assign font[3][99] = 14'b00000000000000;
	assign font[4][99] = 14'b00000000000000;
	assign font[5][99] = 14'b00000000000000;
	assign font[6][99] = 14'b00000000000000;
	assign font[7][99] = 14'b00000000000000;
	assign font[8][99] = 14'b00000000000000;
	assign font[9][99] = 14'b00000000000000;
	assign font[10][99] = 14'b00000000000000;
	assign font[11][99] = 14'b00000000000000;
	assign font[12][99] = 14'b00000000000000;
	assign font[13][99] = 14'b00000000000000;
	assign font[14][99] = 14'b00000111111000;
	assign font[15][99] = 14'b00000111111000;
	assign font[16][99] = 14'b00000100001000;
	assign font[17][99] = 14'b00011100001110;
	assign font[18][99] = 14'b00011100001110;
	assign font[19][99] = 14'b00111000000000;
	assign font[20][99] = 14'b00111000000000;
	assign font[21][99] = 14'b00111000000000;
	assign font[22][99] = 14'b00011100001110;
	assign font[23][99] = 14'b00011100001110;
	assign font[24][99] = 14'b00000100001000;
	assign font[25][99] = 14'b00000111111000;
	assign font[26][99] = 14'b00000111111000;
	assign font[27][99] = 14'b00000000000000;
	assign font[28][99] = 14'b00000000000000;
	assign font[29][99] = 14'b00000000000000;
	assign font[30][99] = 14'b00000000000000;
	assign font[31][99] = 14'b00000000000000;

	assign font[0][100] = 14'b00000000000000;
	assign font[1][100] = 14'b00000000000000;
	assign font[2][100] = 14'b00000000000000;
	assign font[3][100] = 14'b00000000000000;
	assign font[4][100] = 14'b00000000000000;
	assign font[5][100] = 14'b00000000000000;
	assign font[6][100] = 14'b00000000000000;
	assign font[7][100] = 14'b00000000000000;
	assign font[8][100] = 14'b00000000000000;
	assign font[9][100] = 14'b00000000001110;
	assign font[10][100] = 14'b00000000001110;
	assign font[11][100] = 14'b00000000001110;
	assign font[12][100] = 14'b00000000001110;
	assign font[13][100] = 14'b00000000001110;
	assign font[14][100] = 14'b00000111111110;
	assign font[15][100] = 14'b00000111111110;
	assign font[16][100] = 14'b00011100001110;
	assign font[17][100] = 14'b00011100001110;
	assign font[18][100] = 14'b00011100001110;
	assign font[19][100] = 14'b00111000001110;
	assign font[20][100] = 14'b00111000001110;
	assign font[21][100] = 14'b00111000001110;
	assign font[22][100] = 14'b00011100001110;
	assign font[23][100] = 14'b00011100001110;
	assign font[24][100] = 14'b00011100001110;
	assign font[25][100] = 14'b00000111111110;
	assign font[26][100] = 14'b00000111111110;
	assign font[27][100] = 14'b00000000000000;
	assign font[28][100] = 14'b00000000000000;
	assign font[29][100] = 14'b00000000000000;
	assign font[30][100] = 14'b00000000000000;
	assign font[31][100] = 14'b00000000000000;

	assign font[0][101] = 14'b00000000000000;
	assign font[1][101] = 14'b00000000000000;
	assign font[2][101] = 14'b00000000000000;
	assign font[3][101] = 14'b00000000000000;
	assign font[4][101] = 14'b00000000000000;
	assign font[5][101] = 14'b00000000000000;
	assign font[6][101] = 14'b00000000000000;
	assign font[7][101] = 14'b00000000000000;
	assign font[8][101] = 14'b00000000000000;
	assign font[9][101] = 14'b00000000000000;
	assign font[10][101] = 14'b00000000000000;
	assign font[11][101] = 14'b00000000000000;
	assign font[12][101] = 14'b00000000000000;
	assign font[13][101] = 14'b00000000000000;
	assign font[14][101] = 14'b00000111111000;
	assign font[15][101] = 14'b00000111111000;
	assign font[16][101] = 14'b00000111111000;
	assign font[17][101] = 14'b00011100001110;
	assign font[18][101] = 14'b00011100001110;
	assign font[19][101] = 14'b00111111111110;
	assign font[20][101] = 14'b00111111111110;
	assign font[21][101] = 14'b00111111111110;
	assign font[22][101] = 14'b00011100000000;
	assign font[23][101] = 14'b00011100000000;
	assign font[24][101] = 14'b00011100000000;
	assign font[25][101] = 14'b00000111111100;
	assign font[26][101] = 14'b00000111111100;
	assign font[27][101] = 14'b00000000000000;
	assign font[28][101] = 14'b00000000000000;
	assign font[29][101] = 14'b00000000000000;
	assign font[30][101] = 14'b00000000000000;
	assign font[31][101] = 14'b00000000000000;

	assign font[0][102] = 14'b00000000000000;
	assign font[1][102] = 14'b00000000000000;
	assign font[2][102] = 14'b00000000000000;
	assign font[3][102] = 14'b00000000000000;
	assign font[4][102] = 14'b00000000000000;
	assign font[5][102] = 14'b00000000000000;
	assign font[6][102] = 14'b00000000000000;
	assign font[7][102] = 14'b00000000000000;
	assign font[8][102] = 14'b00000000000000;
	assign font[9][102] = 14'b00000111111000;
	assign font[10][102] = 14'b00000111111000;
	assign font[11][102] = 14'b00001110000000;
	assign font[12][102] = 14'b00001110000000;
	assign font[13][102] = 14'b00001110000000;
	assign font[14][102] = 14'b00111111111000;
	assign font[15][102] = 14'b00111111111000;
	assign font[16][102] = 14'b00111111111000;
	assign font[17][102] = 14'b00001110000000;
	assign font[18][102] = 14'b00001110000000;
	assign font[19][102] = 14'b00001110000000;
	assign font[20][102] = 14'b00001110000000;
	assign font[21][102] = 14'b00001110000000;
	assign font[22][102] = 14'b00001110000000;
	assign font[23][102] = 14'b00001110000000;
	assign font[24][102] = 14'b00001110000000;
	assign font[25][102] = 14'b00011111100000;
	assign font[26][102] = 14'b00011111100000;
	assign font[27][102] = 14'b00000000000000;
	assign font[28][102] = 14'b00000000000000;
	assign font[29][102] = 14'b00000000000000;
	assign font[30][102] = 14'b00000000000000;
	assign font[31][102] = 14'b00000000000000;

	assign font[0][103] = 14'b00000000000000;
	assign font[1][103] = 14'b00000000000000;
	assign font[2][103] = 14'b00000000000000;
	assign font[3][103] = 14'b00000000000000;
	assign font[4][103] = 14'b00000000000000;
	assign font[5][103] = 14'b00000000000000;
	assign font[6][103] = 14'b00000000000000;
	assign font[7][103] = 14'b00000000000000;
	assign font[8][103] = 14'b00000000000000;
	assign font[9][103] = 14'b00000000000000;
	assign font[10][103] = 14'b00000000000000;
	assign font[11][103] = 14'b00000000000000;
	assign font[12][103] = 14'b00000000000000;
	assign font[13][103] = 14'b00000000000000;
	assign font[14][103] = 14'b00000111111110;
	assign font[15][103] = 14'b00000111111110;
	assign font[16][103] = 14'b00011100001110;
	assign font[17][103] = 14'b00011100001110;
	assign font[18][103] = 14'b00011100001110;
	assign font[19][103] = 14'b00111000001110;
	assign font[20][103] = 14'b00111000001110;
	assign font[21][103] = 14'b00011100001110;
	assign font[22][103] = 14'b00011100001110;
	assign font[23][103] = 14'b00011100001110;
	assign font[24][103] = 14'b00000111111110;
	assign font[25][103] = 14'b00000111111110;
	assign font[26][103] = 14'b00000111111110;
	assign font[27][103] = 14'b00000000001100;
	assign font[28][103] = 14'b00000000001100;
	assign font[29][103] = 14'b00000000001100;
	assign font[30][103] = 14'b00000111111000;
	assign font[31][103] = 14'b00000111111000;

	assign font[0][104] = 14'b00000000000000;
	assign font[1][104] = 14'b00000000000000;
	assign font[2][104] = 14'b00000000000000;
	assign font[3][104] = 14'b00000000000000;
	assign font[4][104] = 14'b00000000000000;
	assign font[5][104] = 14'b00000000000000;
	assign font[6][104] = 14'b00000000000000;
	assign font[7][104] = 14'b00000000000000;
	assign font[8][104] = 14'b00000000000000;
	assign font[9][104] = 14'b00111000000000;
	assign font[10][104] = 14'b00111000000000;
	assign font[11][104] = 14'b00111000000000;
	assign font[12][104] = 14'b00111000000000;
	assign font[13][104] = 14'b00111000000000;
	assign font[14][104] = 14'b00111111111000;
	assign font[15][104] = 14'b00111111111000;
	assign font[16][104] = 14'b00111000001000;
	assign font[17][104] = 14'b00111100001110;
	assign font[18][104] = 14'b00111100001110;
	assign font[19][104] = 14'b00111000001110;
	assign font[20][104] = 14'b00111000001110;
	assign font[21][104] = 14'b00111000001110;
	assign font[22][104] = 14'b00111000001110;
	assign font[23][104] = 14'b00111000001110;
	assign font[24][104] = 14'b00111000001110;
	assign font[25][104] = 14'b00111000001110;
	assign font[26][104] = 14'b00111000001110;
	assign font[27][104] = 14'b00000000000000;
	assign font[28][104] = 14'b00000000000000;
	assign font[29][104] = 14'b00000000000000;
	assign font[30][104] = 14'b00000000000000;
	assign font[31][104] = 14'b00000000000000;

	assign font[0][105] = 14'b00000000000000;
	assign font[1][105] = 14'b00000000000000;
	assign font[2][105] = 14'b00000000000000;
	assign font[3][105] = 14'b00000000000000;
	assign font[4][105] = 14'b00000000000000;
	assign font[5][105] = 14'b00000000000000;
	assign font[6][105] = 14'b00000000000000;
	assign font[7][105] = 14'b00000000000000;
	assign font[8][105] = 14'b00000000000000;
	assign font[9][105] = 14'b00000011100000;
	assign font[10][105] = 14'b00000011100000;
	assign font[11][105] = 14'b00000000000000;
	assign font[12][105] = 14'b00000000000000;
	assign font[13][105] = 14'b00000000000000;
	assign font[14][105] = 14'b00001111100000;
	assign font[15][105] = 14'b00001111100000;
	assign font[16][105] = 14'b00000011100000;
	assign font[17][105] = 14'b00000011100000;
	assign font[18][105] = 14'b00000011100000;
	assign font[19][105] = 14'b00000011100000;
	assign font[20][105] = 14'b00000011100000;
	assign font[21][105] = 14'b00000011100000;
	assign font[22][105] = 14'b00000011100000;
	assign font[23][105] = 14'b00000011100000;
	assign font[24][105] = 14'b00000011100000;
	assign font[25][105] = 14'b00011111111000;
	assign font[26][105] = 14'b00011111111000;
	assign font[27][105] = 14'b00000000000000;
	assign font[28][105] = 14'b00000000000000;
	assign font[29][105] = 14'b00000000000000;
	assign font[30][105] = 14'b00000000000000;
	assign font[31][105] = 14'b00000000000000;

	assign font[0][106] = 14'b00000000000000;
	assign font[1][106] = 14'b00000000000000;
	assign font[2][106] = 14'b00000000000000;
	assign font[3][106] = 14'b00000000000000;
	assign font[4][106] = 14'b00000000000000;
	assign font[5][106] = 14'b00000000000000;
	assign font[6][106] = 14'b00000000000000;
	assign font[7][106] = 14'b00000000000000;
	assign font[8][106] = 14'b00000000000000;
	assign font[9][106] = 14'b00000011100000;
	assign font[10][106] = 14'b00000011100000;
	assign font[11][106] = 14'b00000000000000;
	assign font[12][106] = 14'b00000000000000;
	assign font[13][106] = 14'b00000000000000;
	assign font[14][106] = 14'b00001111100000;
	assign font[15][106] = 14'b00001111100000;
	assign font[16][106] = 14'b00000011100000;
	assign font[17][106] = 14'b00000011100000;
	assign font[18][106] = 14'b00000011100000;
	assign font[19][106] = 14'b00000011100000;
	assign font[20][106] = 14'b00000011100000;
	assign font[21][106] = 14'b00000011100000;
	assign font[22][106] = 14'b00000011100000;
	assign font[23][106] = 14'b00000011100000;
	assign font[24][106] = 14'b00000011100000;
	assign font[25][106] = 14'b00000011100000;
	assign font[26][106] = 14'b00000011100000;
	assign font[27][106] = 14'b00000111100000;
	assign font[28][106] = 14'b00000111100000;
	assign font[29][106] = 14'b00000111100000;
	assign font[30][106] = 14'b00111111000000;
	assign font[31][106] = 14'b00111111000000;

	assign font[0][107] = 14'b00000000000000;
	assign font[1][107] = 14'b00000000000000;
	assign font[2][107] = 14'b00000000000000;
	assign font[3][107] = 14'b00000000000000;
	assign font[4][107] = 14'b00000000000000;
	assign font[5][107] = 14'b00000000000000;
	assign font[6][107] = 14'b00000000000000;
	assign font[7][107] = 14'b00000000000000;
	assign font[8][107] = 14'b00000000000000;
	assign font[9][107] = 14'b00111000000000;
	assign font[10][107] = 14'b00111000000000;
	assign font[11][107] = 14'b00111000000000;
	assign font[12][107] = 14'b00111000000000;
	assign font[13][107] = 14'b00111000000000;
	assign font[14][107] = 14'b00111000111100;
	assign font[15][107] = 14'b00111000111100;
	assign font[16][107] = 14'b00111011100000;
	assign font[17][107] = 14'b00111011100000;
	assign font[18][107] = 14'b00111011100000;
	assign font[19][107] = 14'b00111111000000;
	assign font[20][107] = 14'b00111111000000;
	assign font[21][107] = 14'b00111011110000;
	assign font[22][107] = 14'b00111011110000;
	assign font[23][107] = 14'b00111011110000;
	assign font[24][107] = 14'b00111011110000;
	assign font[25][107] = 14'b00111000111110;
	assign font[26][107] = 14'b00111000111110;
	assign font[27][107] = 14'b00000000000000;
	assign font[28][107] = 14'b00000000000000;
	assign font[29][107] = 14'b00000000000000;
	assign font[30][107] = 14'b00000000000000;
	assign font[31][107] = 14'b00000000000000;

	assign font[0][108] = 14'b00000000000000;
	assign font[1][108] = 14'b00000000000000;
	assign font[2][108] = 14'b00000000000000;
	assign font[3][108] = 14'b00000000000000;
	assign font[4][108] = 14'b00000000000000;
	assign font[5][108] = 14'b00000000000000;
	assign font[6][108] = 14'b00000000000000;
	assign font[7][108] = 14'b00000000000000;
	assign font[8][108] = 14'b00000000000000;
	assign font[9][108] = 14'b00001111100000;
	assign font[10][108] = 14'b00001111100000;
	assign font[11][108] = 14'b00000011100000;
	assign font[12][108] = 14'b00000011100000;
	assign font[13][108] = 14'b00000011100000;
	assign font[14][108] = 14'b00000011100000;
	assign font[15][108] = 14'b00000011100000;
	assign font[16][108] = 14'b00000011100000;
	assign font[17][108] = 14'b00000011100000;
	assign font[18][108] = 14'b00000011100000;
	assign font[19][108] = 14'b00000011100000;
	assign font[20][108] = 14'b00000011100000;
	assign font[21][108] = 14'b00000011100000;
	assign font[22][108] = 14'b00000011100000;
	assign font[23][108] = 14'b00000011100000;
	assign font[24][108] = 14'b00000011100000;
	assign font[25][108] = 14'b00011111111100;
	assign font[26][108] = 14'b00001111111100;
	assign font[27][108] = 14'b00000000000000;
	assign font[28][108] = 14'b00000000000000;
	assign font[29][108] = 14'b00000000000000;
	assign font[30][108] = 14'b00000000000000;
	assign font[31][108] = 14'b00000000000000;

	assign font[0][109] = 14'b00000000000000;
	assign font[1][109] = 14'b00000000000000;
	assign font[2][109] = 14'b00000000000000;
	assign font[3][109] = 14'b00000000000000;
	assign font[4][109] = 14'b00000000000000;
	assign font[5][109] = 14'b00000000000000;
	assign font[6][109] = 14'b00000000000000;
	assign font[7][109] = 14'b00000000000000;
	assign font[8][109] = 14'b00000000000000;
	assign font[9][109] = 14'b00000000000000;
	assign font[10][109] = 14'b00000000000000;
	assign font[11][109] = 14'b00000000000000;
	assign font[12][109] = 14'b00000000000000;
	assign font[13][109] = 14'b00000000000000;
	assign font[14][109] = 14'b00110111111100;
	assign font[15][109] = 14'b00110111111100;
	assign font[16][109] = 14'b00111011001110;
	assign font[17][109] = 14'b00111011001110;
	assign font[18][109] = 14'b00111011001110;
	assign font[19][109] = 14'b00111011001110;
	assign font[20][109] = 14'b00111011001110;
	assign font[21][109] = 14'b00111011001110;
	assign font[22][109] = 14'b00111011001110;
	assign font[23][109] = 14'b00111011001110;
	assign font[24][109] = 14'b00111011001110;
	assign font[25][109] = 14'b00111011001110;
	assign font[26][109] = 14'b00111011001110;
	assign font[27][109] = 14'b00000000000000;
	assign font[28][109] = 14'b00000000000000;
	assign font[29][109] = 14'b00000000000000;
	assign font[30][109] = 14'b00000000000000;
	assign font[31][109] = 14'b00000000000000;

	assign font[0][110] = 14'b00000000000000;
	assign font[1][110] = 14'b00000000000000;
	assign font[2][110] = 14'b00000000000000;
	assign font[3][110] = 14'b00000000000000;
	assign font[4][110] = 14'b00000000000000;
	assign font[5][110] = 14'b00000000000000;
	assign font[6][110] = 14'b00000000000000;
	assign font[7][110] = 14'b00000000000000;
	assign font[8][110] = 14'b00000000000000;
	assign font[9][110] = 14'b00000000000000;
	assign font[10][110] = 14'b00000000000000;
	assign font[11][110] = 14'b00000000000000;
	assign font[12][110] = 14'b00000000000000;
	assign font[13][110] = 14'b00000000000000;
	assign font[14][110] = 14'b00111111111000;
	assign font[15][110] = 14'b00111111111000;
	assign font[16][110] = 14'b00111000001000;
	assign font[17][110] = 14'b00111100001110;
	assign font[18][110] = 14'b00111100001110;
	assign font[19][110] = 14'b00111000001110;
	assign font[20][110] = 14'b00111000001110;
	assign font[21][110] = 14'b00111000001110;
	assign font[22][110] = 14'b00111000001110;
	assign font[23][110] = 14'b00111000001110;
	assign font[24][110] = 14'b00111000001110;
	assign font[25][110] = 14'b00111000001110;
	assign font[26][110] = 14'b00111000001110;
	assign font[27][110] = 14'b00000000000000;
	assign font[28][110] = 14'b00000000000000;
	assign font[29][110] = 14'b00000000000000;
	assign font[30][110] = 14'b00000000000000;
	assign font[31][110] = 14'b00000000000000;

	assign font[0][111] = 14'b00000000000000;
	assign font[1][111] = 14'b00000000000000;
	assign font[2][111] = 14'b00000000000000;
	assign font[3][111] = 14'b00000000000000;
	assign font[4][111] = 14'b00000000000000;
	assign font[5][111] = 14'b00000000000000;
	assign font[6][111] = 14'b00000000000000;
	assign font[7][111] = 14'b00000000000000;
	assign font[8][111] = 14'b00000000000000;
	assign font[9][111] = 14'b00000000000000;
	assign font[10][111] = 14'b00000000000000;
	assign font[11][111] = 14'b00000000000000;
	assign font[12][111] = 14'b00000000000000;
	assign font[13][111] = 14'b00000000000000;
	assign font[14][111] = 14'b00000111111000;
	assign font[15][111] = 14'b00000111111000;
	assign font[16][111] = 14'b00011100011100;
	assign font[17][111] = 14'b00011100011100;
	assign font[18][111] = 14'b00011100011100;
	assign font[19][111] = 14'b00111000001110;
	assign font[20][111] = 14'b00111000001110;
	assign font[21][111] = 14'b00011100011100;
	assign font[22][111] = 14'b00011100011100;
	assign font[23][111] = 14'b00011100011100;
	assign font[24][111] = 14'b00000100011000;
	assign font[25][111] = 14'b00000111111000;
	assign font[26][111] = 14'b00000111111000;
	assign font[27][111] = 14'b00000000000000;
	assign font[28][111] = 14'b00000000000000;
	assign font[29][111] = 14'b00000000000000;
	assign font[30][111] = 14'b00000000000000;
	assign font[31][111] = 14'b00000000000000;

	assign font[0][112] = 14'b00000000000000;
	assign font[1][112] = 14'b00000000000000;
	assign font[2][112] = 14'b00000000000000;
	assign font[3][112] = 14'b00000000000000;
	assign font[4][112] = 14'b00000000000000;
	assign font[5][112] = 14'b00000000000000;
	assign font[6][112] = 14'b00000000000000;
	assign font[7][112] = 14'b00000000000000;
	assign font[8][112] = 14'b00000000000000;
	assign font[9][112] = 14'b00000000000000;
	assign font[10][112] = 14'b00000000000000;
	assign font[11][112] = 14'b00000000000000;
	assign font[12][112] = 14'b00000000000000;
	assign font[13][112] = 14'b00000000000000;
	assign font[14][112] = 14'b00111111110000;
	assign font[15][112] = 14'b00111111110000;
	assign font[16][112] = 14'b00111100011100;
	assign font[17][112] = 14'b00111100011100;
	assign font[18][112] = 14'b00111100011100;
	assign font[19][112] = 14'b00111000001110;
	assign font[20][112] = 14'b00111000001110;
	assign font[21][112] = 14'b00111000011100;
	assign font[22][112] = 14'b00111000011100;
	assign font[23][112] = 14'b00111000011100;
	assign font[24][112] = 14'b00111000010000;
	assign font[25][112] = 14'b00111111110000;
	assign font[26][112] = 14'b00111111110000;
	assign font[27][112] = 14'b00111000000000;
	assign font[28][112] = 14'b00111000000000;
	assign font[29][112] = 14'b00111000000000;
	assign font[30][112] = 14'b00111000000000;
	assign font[31][112] = 14'b00111000000000;

	assign font[0][113] = 14'b00000000000000;
	assign font[1][113] = 14'b00000000000000;
	assign font[2][113] = 14'b00000000000000;
	assign font[3][113] = 14'b00000000000000;
	assign font[4][113] = 14'b00000000000000;
	assign font[5][113] = 14'b00000000000000;
	assign font[6][113] = 14'b00000000000000;
	assign font[7][113] = 14'b00000000000000;
	assign font[8][113] = 14'b00000000000000;
	assign font[9][113] = 14'b00000000000000;
	assign font[10][113] = 14'b00000000000000;
	assign font[11][113] = 14'b00000000000000;
	assign font[12][113] = 14'b00000000000000;
	assign font[13][113] = 14'b00000000000000;
	assign font[14][113] = 14'b00000111111110;
	assign font[15][113] = 14'b00000111111110;
	assign font[16][113] = 14'b00011100001110;
	assign font[17][113] = 14'b00011100001110;
	assign font[18][113] = 14'b00011100001110;
	assign font[19][113] = 14'b00111000001110;
	assign font[20][113] = 14'b00111000001110;
	assign font[21][113] = 14'b00111000001110;
	assign font[22][113] = 14'b00011100001110;
	assign font[23][113] = 14'b00011100001110;
	assign font[24][113] = 14'b00011100001110;
	assign font[25][113] = 14'b00000111111110;
	assign font[26][113] = 14'b00000111111110;
	assign font[27][113] = 14'b00000000001110;
	assign font[28][113] = 14'b00000000001110;
	assign font[29][113] = 14'b00000000001110;
	assign font[30][113] = 14'b00000000001110;
	assign font[31][113] = 14'b00000000001110;

	assign font[0][114] = 14'b00000000000000;
	assign font[1][114] = 14'b00000000000000;
	assign font[2][114] = 14'b00000000000000;
	assign font[3][114] = 14'b00000000000000;
	assign font[4][114] = 14'b00000000000000;
	assign font[5][114] = 14'b00000000000000;
	assign font[6][114] = 14'b00000000000000;
	assign font[7][114] = 14'b00000000000000;
	assign font[8][114] = 14'b00000000000000;
	assign font[9][114] = 14'b00000000000000;
	assign font[10][114] = 14'b00000000000000;
	assign font[11][114] = 14'b00000000000000;
	assign font[12][114] = 14'b00000000000000;
	assign font[13][114] = 14'b00000000000000;
	assign font[14][114] = 14'b00111111111100;
	assign font[15][114] = 14'b00111111111100;
	assign font[16][114] = 14'b00001111001110;
	assign font[17][114] = 14'b00001111001110;
	assign font[18][114] = 14'b00001111001110;
	assign font[19][114] = 14'b00001110000000;
	assign font[20][114] = 14'b00001110000000;
	assign font[21][114] = 14'b00001110000000;
	assign font[22][114] = 14'b00001110000000;
	assign font[23][114] = 14'b00001110000000;
	assign font[24][114] = 14'b00001110000000;
	assign font[25][114] = 14'b00111111100000;
	assign font[26][114] = 14'b00111111100000;
	assign font[27][114] = 14'b00000000000000;
	assign font[28][114] = 14'b00000000000000;
	assign font[29][114] = 14'b00000000000000;
	assign font[30][114] = 14'b00000000000000;
	assign font[31][114] = 14'b00000000000000;

	assign font[0][115] = 14'b00000000000000;
	assign font[1][115] = 14'b00000000000000;
	assign font[2][115] = 14'b00000000000000;
	assign font[3][115] = 14'b00000000000000;
	assign font[4][115] = 14'b00000000000000;
	assign font[5][115] = 14'b00000000000000;
	assign font[6][115] = 14'b00000000000000;
	assign font[7][115] = 14'b00000000000000;
	assign font[8][115] = 14'b00000000000000;
	assign font[9][115] = 14'b00000000000000;
	assign font[10][115] = 14'b00000000000000;
	assign font[11][115] = 14'b00000000000000;
	assign font[12][115] = 14'b00000000000000;
	assign font[13][115] = 14'b00000000000000;
	assign font[14][115] = 14'b00001111111000;
	assign font[15][115] = 14'b00001111111000;
	assign font[16][115] = 14'b00111000000000;
	assign font[17][115] = 14'b00111000000000;
	assign font[18][115] = 14'b00111000000000;
	assign font[19][115] = 14'b00001111110000;
	assign font[20][115] = 14'b00001111110000;
	assign font[21][115] = 14'b00001111110000;
	assign font[22][115] = 14'b00000000011100;
	assign font[23][115] = 14'b00000000011100;
	assign font[24][115] = 14'b00000000010000;
	assign font[25][115] = 14'b00011111110000;
	assign font[26][115] = 14'b00011111110000;
	assign font[27][115] = 14'b00000000000000;
	assign font[28][115] = 14'b00000000000000;
	assign font[29][115] = 14'b00000000000000;
	assign font[30][115] = 14'b00000000000000;
	assign font[31][115] = 14'b00000000000000;

	assign font[0][116] = 14'b00000000000000;
	assign font[1][116] = 14'b00000000000000;
	assign font[2][116] = 14'b00000000000000;
	assign font[3][116] = 14'b00000000000000;
	assign font[4][116] = 14'b00000000000000;
	assign font[5][116] = 14'b00000000000000;
	assign font[6][116] = 14'b00000000000000;
	assign font[7][116] = 14'b00000000000000;
	assign font[8][116] = 14'b00000000000000;
	assign font[9][116] = 14'b00000111000000;
	assign font[10][116] = 14'b00000111000000;
	assign font[11][116] = 14'b00000111000000;
	assign font[12][116] = 14'b00000111000000;
	assign font[13][116] = 14'b00000111000000;
	assign font[14][116] = 14'b00111111111000;
	assign font[15][116] = 14'b00111111111000;
	assign font[16][116] = 14'b00000111000000;
	assign font[17][116] = 14'b00000111000000;
	assign font[18][116] = 14'b00000111000000;
	assign font[19][116] = 14'b00000111000000;
	assign font[20][116] = 14'b00000111000000;
	assign font[21][116] = 14'b00000111000000;
	assign font[22][116] = 14'b00000111000000;
	assign font[23][116] = 14'b00000111000000;
	assign font[24][116] = 14'b00000111000000;
	assign font[25][116] = 14'b00000111111000;
	assign font[26][116] = 14'b00000111111000;
	assign font[27][116] = 14'b00000000000000;
	assign font[28][116] = 14'b00000000000000;
	assign font[29][116] = 14'b00000000000000;
	assign font[30][116] = 14'b00000000000000;
	assign font[31][116] = 14'b00000000000000;

	assign font[0][117] = 14'b00000000000000;
	assign font[1][117] = 14'b00000000000000;
	assign font[2][117] = 14'b00000000000000;
	assign font[3][117] = 14'b00000000000000;
	assign font[4][117] = 14'b00000000000000;
	assign font[5][117] = 14'b00000000000000;
	assign font[6][117] = 14'b00000000000000;
	assign font[7][117] = 14'b00000000000000;
	assign font[8][117] = 14'b00000000000000;
	assign font[9][117] = 14'b00000000000000;
	assign font[10][117] = 14'b00000000000000;
	assign font[11][117] = 14'b00000000000000;
	assign font[12][117] = 14'b00000000000000;
	assign font[13][117] = 14'b00000000000000;
	assign font[14][117] = 14'b00111000001110;
	assign font[15][117] = 14'b00111000001110;
	assign font[16][117] = 14'b00111000001110;
	assign font[17][117] = 14'b00111000001110;
	assign font[18][117] = 14'b00111000001110;
	assign font[19][117] = 14'b00111000001110;
	assign font[20][117] = 14'b00111000001110;
	assign font[21][117] = 14'b00111100001110;
	assign font[22][117] = 14'b00111100001110;
	assign font[23][117] = 14'b00111100001110;
	assign font[24][117] = 14'b00001100001110;
	assign font[25][117] = 14'b00001111111110;
	assign font[26][117] = 14'b00001111111110;
	assign font[27][117] = 14'b00000000000000;
	assign font[28][117] = 14'b00000000000000;
	assign font[29][117] = 14'b00000000000000;
	assign font[30][117] = 14'b00000000000000;
	assign font[31][117] = 14'b00000000000000;

	assign font[0][118] = 14'b00000000000000;
	assign font[1][118] = 14'b00000000000000;
	assign font[2][118] = 14'b00000000000000;
	assign font[3][118] = 14'b00000000000000;
	assign font[4][118] = 14'b00000000000000;
	assign font[5][118] = 14'b00000000000000;
	assign font[6][118] = 14'b00000000000000;
	assign font[7][118] = 14'b00000000000000;
	assign font[8][118] = 14'b00000000000000;
	assign font[9][118] = 14'b00000000000000;
	assign font[10][118] = 14'b00000000000000;
	assign font[11][118] = 14'b00000000000000;
	assign font[12][118] = 14'b00000000000000;
	assign font[13][118] = 14'b00000000000000;
	assign font[14][118] = 14'b00111000011100;
	assign font[15][118] = 14'b00111000011100;
	assign font[16][118] = 14'b00111000011100;
	assign font[17][118] = 14'b00011100011000;
	assign font[18][118] = 14'b00011100011000;
	assign font[19][118] = 14'b00001110111000;
	assign font[20][118] = 14'b00001110111000;
	assign font[21][118] = 14'b00001110111000;
	assign font[22][118] = 14'b00000111110000;
	assign font[23][118] = 14'b00000111110000;
	assign font[24][118] = 14'b00000111110000;
	assign font[25][118] = 14'b00000011100000;
	assign font[26][118] = 14'b00000011100000;
	assign font[27][118] = 14'b00000000000000;
	assign font[28][118] = 14'b00000000000000;
	assign font[29][118] = 14'b00000000000000;
	assign font[30][118] = 14'b00000000000000;
	assign font[31][118] = 14'b00000000000000;

	assign font[0][119] = 14'b00000000000000;
	assign font[1][119] = 14'b00000000000000;
	assign font[2][119] = 14'b00000000000000;
	assign font[3][119] = 14'b00000000000000;
	assign font[4][119] = 14'b00000000000000;
	assign font[5][119] = 14'b00000000000000;
	assign font[6][119] = 14'b00000000000000;
	assign font[7][119] = 14'b00000000000000;
	assign font[8][119] = 14'b00000000000000;
	assign font[9][119] = 14'b00000000000000;
	assign font[10][119] = 14'b00000000000000;
	assign font[11][119] = 14'b00000000000000;
	assign font[12][119] = 14'b00000000000000;
	assign font[13][119] = 14'b00000000000000;
	assign font[14][119] = 14'b00111011001110;
	assign font[15][119] = 14'b00111011001110;
	assign font[16][119] = 14'b00111011001110;
	assign font[17][119] = 14'b00111011001110;
	assign font[18][119] = 14'b00111011001110;
	assign font[19][119] = 14'b00011011101100;
	assign font[20][119] = 14'b00011011101100;
	assign font[21][119] = 14'b00011011101100;
	assign font[22][119] = 14'b00011110111100;
	assign font[23][119] = 14'b00011110111100;
	assign font[24][119] = 14'b00001100011000;
	assign font[25][119] = 14'b00001100011000;
	assign font[26][119] = 14'b00001100011000;
	assign font[27][119] = 14'b00000000000000;
	assign font[28][119] = 14'b00000000000000;
	assign font[29][119] = 14'b00000000000000;
	assign font[30][119] = 14'b00000000000000;
	assign font[31][119] = 14'b00000000000000;

	assign font[0][120] = 14'b00000000000000;
	assign font[1][120] = 14'b00000000000000;
	assign font[2][120] = 14'b00000000000000;
	assign font[3][120] = 14'b00000000000000;
	assign font[4][120] = 14'b00000000000000;
	assign font[5][120] = 14'b00000000000000;
	assign font[6][120] = 14'b00000000000000;
	assign font[7][120] = 14'b00000000000000;
	assign font[8][120] = 14'b00000000000000;
	assign font[9][120] = 14'b00000000000000;
	assign font[10][120] = 14'b00000000000000;
	assign font[11][120] = 14'b00000000000000;
	assign font[12][120] = 14'b00000000000000;
	assign font[13][120] = 14'b00000000000000;
	assign font[14][120] = 14'b00011100011100;
	assign font[15][120] = 14'b00011100011100;
	assign font[16][120] = 14'b00001110111000;
	assign font[17][120] = 14'b00001110111000;
	assign font[18][120] = 14'b00001110111000;
	assign font[19][120] = 14'b00000010110000;
	assign font[20][120] = 14'b00000011110000;
	assign font[21][120] = 14'b00000011110000;
	assign font[22][120] = 14'b00001110111000;
	assign font[23][120] = 14'b00001110111000;
	assign font[24][120] = 14'b00001100011100;
	assign font[25][120] = 14'b00011100011100;
	assign font[26][120] = 14'b00011100011100;
	assign font[27][120] = 14'b00000000000000;
	assign font[28][120] = 14'b00000000000000;
	assign font[29][120] = 14'b00000000000000;
	assign font[30][120] = 14'b00000000000000;
	assign font[31][120] = 14'b00000000000000;

	assign font[0][121] = 14'b00000000000000;
	assign font[1][121] = 14'b00000000000000;
	assign font[2][121] = 14'b00000000000000;
	assign font[3][121] = 14'b00000000000000;
	assign font[4][121] = 14'b00000000000000;
	assign font[5][121] = 14'b00000000000000;
	assign font[6][121] = 14'b00000000000000;
	assign font[7][121] = 14'b00000000000000;
	assign font[8][121] = 14'b00000000000000;
	assign font[9][121] = 14'b00000000000000;
	assign font[10][121] = 14'b00000000000000;
	assign font[11][121] = 14'b00000000000000;
	assign font[12][121] = 14'b00000000000000;
	assign font[13][121] = 14'b00000000000000;
	assign font[14][121] = 14'b00111000001110;
	assign font[15][121] = 14'b00111000001110;
	assign font[16][121] = 14'b00011100001100;
	assign font[17][121] = 14'b00011100001100;
	assign font[18][121] = 14'b00011100001100;
	assign font[19][121] = 14'b00001110111000;
	assign font[20][121] = 14'b00001110111000;
	assign font[21][121] = 14'b00001110111000;
	assign font[22][121] = 14'b00000111110000;
	assign font[23][121] = 14'b00000111110000;
	assign font[24][121] = 14'b00000011110000;
	assign font[25][121] = 14'b00000011110000;
	assign font[26][121] = 14'b00000011110000;
	assign font[27][121] = 14'b00000011100000;
	assign font[28][121] = 14'b00000011100000;
	assign font[29][121] = 14'b00000010000000;
	assign font[30][121] = 14'b00011110000000;
	assign font[31][121] = 14'b00011110000000;

	assign font[0][122] = 14'b00000000000000;
	assign font[1][122] = 14'b00000000000000;
	assign font[2][122] = 14'b00000000000000;
	assign font[3][122] = 14'b00000000000000;
	assign font[4][122] = 14'b00000000000000;
	assign font[5][122] = 14'b00000000000000;
	assign font[6][122] = 14'b00000000000000;
	assign font[7][122] = 14'b00000000000000;
	assign font[8][122] = 14'b00000000000000;
	assign font[9][122] = 14'b00000000000000;
	assign font[10][122] = 14'b00000000000000;
	assign font[11][122] = 14'b00000000000000;
	assign font[12][122] = 14'b00000000000000;
	assign font[13][122] = 14'b00000000000000;
	assign font[14][122] = 14'b00111111111000;
	assign font[15][122] = 14'b00111111111000;
	assign font[16][122] = 14'b00000001110000;
	assign font[17][122] = 14'b00000001110000;
	assign font[18][122] = 14'b00000001110000;
	assign font[19][122] = 14'b00000111000000;
	assign font[20][122] = 14'b00000111000000;
	assign font[21][122] = 14'b00000111000000;
	assign font[22][122] = 14'b00111000000000;
	assign font[23][122] = 14'b00111000000000;
	assign font[24][122] = 14'b00111000000000;
	assign font[25][122] = 14'b00111111111000;
	assign font[26][122] = 14'b00111111111000;
	assign font[27][122] = 14'b00000000000000;
	assign font[28][122] = 14'b00000000000000;
	assign font[29][122] = 14'b00000000000000;
	assign font[30][122] = 14'b00000000000000;
	assign font[31][122] = 14'b00000000000000;

	assign font[0][123] = 14'b00000000000000;
	assign font[1][123] = 14'b00000000000000;
	assign font[2][123] = 14'b00000000000000;
	assign font[3][123] = 14'b00000000000000;
	assign font[4][123] = 14'b00000000000000;
	assign font[5][123] = 14'b00000000000000;
	assign font[6][123] = 14'b00000000111100;
	assign font[7][123] = 14'b00000000111100;
	assign font[8][123] = 14'b00000000110000;
	assign font[9][123] = 14'b00000001110000;
	assign font[10][123] = 14'b00000001110000;
	assign font[11][123] = 14'b00000011000000;
	assign font[12][123] = 14'b00000011000000;
	assign font[13][123] = 14'b00000011000000;
	assign font[14][123] = 14'b00000011000000;
	assign font[15][123] = 14'b00000011000000;
	assign font[16][123] = 14'b00000000000000;
	assign font[17][123] = 14'b00011100000000;
	assign font[18][123] = 14'b00011100000000;
	assign font[19][123] = 14'b00000011000000;
	assign font[20][123] = 14'b00000011000000;
	assign font[21][123] = 14'b00000011000000;
	assign font[22][123] = 14'b00000011000000;
	assign font[23][123] = 14'b00000011000000;
	assign font[24][123] = 14'b00000001100000;
	assign font[25][123] = 14'b00000001110000;
	assign font[26][123] = 14'b00000001110000;
	assign font[27][123] = 14'b00000000111000;
	assign font[28][123] = 14'b00000000111000;
	assign font[29][123] = 14'b00000000000000;
	assign font[30][123] = 14'b00000000000000;
	assign font[31][123] = 14'b00000000000000;

	assign font[0][124] = 14'b00000000000000;
	assign font[1][124] = 14'b00000000000000;
	assign font[2][124] = 14'b00000000000000;
	assign font[3][124] = 14'b00000000000000;
	assign font[4][124] = 14'b00000000000000;
	assign font[5][124] = 14'b00000000000000;
	assign font[6][124] = 14'b00000000000000;
	assign font[7][124] = 14'b00000011100000;
	assign font[8][124] = 14'b00000011100000;
	assign font[9][124] = 14'b00000011100000;
	assign font[10][124] = 14'b00000011100000;
	assign font[11][124] = 14'b00000011100000;
	assign font[12][124] = 14'b00000011100000;
	assign font[13][124] = 14'b00000011100000;
	assign font[14][124] = 14'b00000011100000;
	assign font[15][124] = 14'b00000011100000;
	assign font[16][124] = 14'b00000011100000;
	assign font[17][124] = 14'b00000011100000;
	assign font[18][124] = 14'b00000011100000;
	assign font[19][124] = 14'b00000011100000;
	assign font[20][124] = 14'b00000011100000;
	assign font[21][124] = 14'b00000011100000;
	assign font[22][124] = 14'b00000011100000;
	assign font[23][124] = 14'b00000011100000;
	assign font[24][124] = 14'b00000011100000;
	assign font[25][124] = 14'b00000011100000;
	assign font[26][124] = 14'b00000011100000;
	assign font[27][124] = 14'b00000011100000;
	assign font[28][124] = 14'b00000011100000;
	assign font[29][124] = 14'b00000011100000;
	assign font[30][124] = 14'b00000000000000;
	assign font[31][124] = 14'b00000000000000;

	assign font[0][125] = 14'b00000000000000;
	assign font[1][125] = 14'b00000000000000;
	assign font[2][125] = 14'b00000000000000;
	assign font[3][125] = 14'b00000000000000;
	assign font[4][125] = 14'b00000000000000;
	assign font[5][125] = 14'b00000000000000;
	assign font[6][125] = 14'b00111000000000;
	assign font[7][125] = 14'b00111000000000;
	assign font[8][125] = 14'b00111000000000;
	assign font[9][125] = 14'b00001110000000;
	assign font[10][125] = 14'b00001110000000;
	assign font[11][125] = 14'b00000011000000;
	assign font[12][125] = 14'b00000011000000;
	assign font[13][125] = 14'b00000011000000;
	assign font[14][125] = 14'b00000011000000;
	assign font[15][125] = 14'b00000011000000;
	assign font[16][125] = 14'b00000011000000;
	assign font[17][125] = 14'b00000000111000;
	assign font[18][125] = 14'b00000000111000;
	assign font[19][125] = 14'b00000011000000;
	assign font[20][125] = 14'b00000011000000;
	assign font[21][125] = 14'b00000011000000;
	assign font[22][125] = 14'b00000011000000;
	assign font[23][125] = 14'b00000011000000;
	assign font[24][125] = 14'b00000010000000;
	assign font[25][125] = 14'b00001110000000;
	assign font[26][125] = 14'b00001110000000;
	assign font[27][125] = 14'b00111000000000;
	assign font[28][125] = 14'b00111000000000;
	assign font[29][125] = 14'b00000000000000;
	assign font[30][125] = 14'b00000000000000;
	assign font[31][125] = 14'b00000000000000;

	assign font[0][126] = 14'b00000000000000;
	assign font[1][126] = 14'b00000000000000;
	assign font[2][126] = 14'b00000000000000;
	assign font[3][126] = 14'b00000000000000;
	assign font[4][126] = 14'b00000000000000;
	assign font[5][126] = 14'b00000000000000;
	assign font[6][126] = 14'b00000000000000;
	assign font[7][126] = 14'b00000000000000;
	assign font[8][126] = 14'b00000000000000;
	assign font[9][126] = 14'b00001111001110;
	assign font[10][126] = 14'b00001111001110;
	assign font[11][126] = 14'b00011111101110;
	assign font[12][126] = 14'b00011111101110;
	assign font[13][126] = 14'b00011111101110;
	assign font[14][126] = 14'b00111011111100;
	assign font[15][126] = 14'b00111011111100;
	assign font[16][126] = 14'b00111011111100;
	assign font[17][126] = 14'b00111001111000;
	assign font[18][126] = 14'b00111001111000;
	assign font[19][126] = 14'b00000000000000;
	assign font[20][126] = 14'b00000000000000;
	assign font[21][126] = 14'b00000000000000;
	assign font[22][126] = 14'b00000000000000;
	assign font[23][126] = 14'b00000000000000;
	assign font[24][126] = 14'b00000000000000;
	assign font[25][126] = 14'b00000000000000;
	assign font[26][126] = 14'b00000000000000;
	assign font[27][126] = 14'b00000000000000;
	assign font[28][126] = 14'b00000000000000;
	assign font[29][126] = 14'b00000000000000;
	assign font[30][126] = 14'b00000000000000;
	assign font[31][126] = 14'b00000000000000;

	assign font[0][127] = 14'b11111111111111;
	assign font[1][127] = 14'b11111111111111;
	assign font[2][127] = 14'b11111111111111;
	assign font[3][127] = 14'b11111111111111;
	assign font[4][127] = 14'b11111111111111;
	assign font[5][127] = 14'b11111111111111;
	assign font[6][127] = 14'b11111111111111;
	assign font[7][127] = 14'b11111111111111;
	assign font[8][127] = 14'b11111111111111;
	assign font[9][127] = 14'b11111111111111;
	assign font[10][127] = 14'b11111111111111;
	assign font[11][127] = 14'b11111111111111;
	assign font[12][127] = 14'b11111111111111;
	assign font[13][127] = 14'b11111111111111;
	assign font[14][127] = 14'b11111111111111;
	assign font[15][127] = 14'b11111111111111;
	assign font[16][127] = 14'b11111111111111;
	assign font[17][127] = 14'b11111111111111;
	assign font[18][127] = 14'b11111111111111;
	assign font[19][127] = 14'b11111111111111;
	assign font[20][127] = 14'b11111111111111;
	assign font[21][127] = 14'b11111111111111;
	assign font[22][127] = 14'b11111111111111;
	assign font[23][127] = 14'b11111111111111;
	assign font[24][127] = 14'b11111111111111;
	assign font[25][127] = 14'b11111111111111;
	assign font[26][127] = 14'b11111111111111;
	assign font[27][127] = 14'b11111111111111;
	assign font[28][127] = 14'b11111111111111;
	assign font[29][127] = 14'b11111111111111;
	assign font[30][127] = 14'b11111111111111;
	assign font[31][127] = 14'b11111111111111;

	assign font[0][128] = 14'b11111111111111;
	assign font[1][128] = 14'b11111111111111;
	assign font[2][128] = 14'b11111111111111;
	assign font[3][128] = 14'b11111111111111;
	assign font[4][128] = 14'b11111111111111;
	assign font[5][128] = 14'b11111111111111;
	assign font[6][128] = 14'b11111111111111;
	assign font[7][128] = 14'b11111111111111;
	assign font[8][128] = 14'b11111111111111;
	assign font[9][128] = 14'b11111111111111;
	assign font[10][128] = 14'b11111111111111;
	assign font[11][128] = 14'b11111111111111;
	assign font[12][128] = 14'b11111111111111;
	assign font[13][128] = 14'b11111111111111;
	assign font[14][128] = 14'b11111111111111;
	assign font[15][128] = 14'b11111111111111;
	assign font[16][128] = 14'b11111111111111;
	assign font[17][128] = 14'b11111111111111;
	assign font[18][128] = 14'b11111111111111;
	assign font[19][128] = 14'b11111111111111;
	assign font[20][128] = 14'b11111111111111;
	assign font[21][128] = 14'b11111111111111;
	assign font[22][128] = 14'b11111111111111;
	assign font[23][128] = 14'b11111111111111;
	assign font[24][128] = 14'b11111111111111;
	assign font[25][128] = 14'b11111111111111;
	assign font[26][128] = 14'b11111111111111;
	assign font[27][128] = 14'b11111111111111;
	assign font[28][128] = 14'b11111111111111;
	assign font[29][128] = 14'b11111111111111;
	assign font[30][128] = 14'b11111111111111;
	assign font[31][128] = 14'b11111111111111;

	assign font[0][129] = 14'b11111111111111;
	assign font[1][129] = 14'b11111111111111;
	assign font[2][129] = 14'b11111111111111;
	assign font[3][129] = 14'b11111111111111;
	assign font[4][129] = 14'b11111111111111;
	assign font[5][129] = 14'b11111111111111;
	assign font[6][129] = 14'b11111111111111;
	assign font[7][129] = 14'b11111111111111;
	assign font[8][129] = 14'b11111111111111;
	assign font[9][129] = 14'b11111111111111;
	assign font[10][129] = 14'b11111111111111;
	assign font[11][129] = 14'b11111111111111;
	assign font[12][129] = 14'b11111111111111;
	assign font[13][129] = 14'b11111111111111;
	assign font[14][129] = 14'b11111111111111;
	assign font[15][129] = 14'b11111111111111;
	assign font[16][129] = 14'b11111111111111;
	assign font[17][129] = 14'b11111111111111;
	assign font[18][129] = 14'b11111111111111;
	assign font[19][129] = 14'b11111111111111;
	assign font[20][129] = 14'b11111111111111;
	assign font[21][129] = 14'b11111111111111;
	assign font[22][129] = 14'b11111111111111;
	assign font[23][129] = 14'b11111111111111;
	assign font[24][129] = 14'b11111111111111;
	assign font[25][129] = 14'b11111111111111;
	assign font[26][129] = 14'b11111111111111;
	assign font[27][129] = 14'b11111111111111;
	assign font[28][129] = 14'b11111111111111;
	assign font[29][129] = 14'b11111111111111;
	assign font[30][129] = 14'b11111111111111;
	assign font[31][129] = 14'b11111111111111;

	assign font[0][130] = 14'b11111111111111;
	assign font[1][130] = 14'b11111111111111;
	assign font[2][130] = 14'b11111111111111;
	assign font[3][130] = 14'b11111111111111;
	assign font[4][130] = 14'b11111111111111;
	assign font[5][130] = 14'b11111111111111;
	assign font[6][130] = 14'b11111111111111;
	assign font[7][130] = 14'b11111111111111;
	assign font[8][130] = 14'b11111111111111;
	assign font[9][130] = 14'b11111111111111;
	assign font[10][130] = 14'b11111111111111;
	assign font[11][130] = 14'b11111111111111;
	assign font[12][130] = 14'b11111111111111;
	assign font[13][130] = 14'b11111111111111;
	assign font[14][130] = 14'b11111111111111;
	assign font[15][130] = 14'b11111111111111;
	assign font[16][130] = 14'b11111111111111;
	assign font[17][130] = 14'b11111111111111;
	assign font[18][130] = 14'b11111111111111;
	assign font[19][130] = 14'b11111111111111;
	assign font[20][130] = 14'b11111111111111;
	assign font[21][130] = 14'b11111111111111;
	assign font[22][130] = 14'b11111111111111;
	assign font[23][130] = 14'b11111111111111;
	assign font[24][130] = 14'b11111111111111;
	assign font[25][130] = 14'b11111111111111;
	assign font[26][130] = 14'b11111111111111;
	assign font[27][130] = 14'b11111111111111;
	assign font[28][130] = 14'b11111111111111;
	assign font[29][130] = 14'b11111111111111;
	assign font[30][130] = 14'b11111111111111;
	assign font[31][130] = 14'b11111111111111;

	assign font[0][131] = 14'b11111111111111;
	assign font[1][131] = 14'b11111111111111;
	assign font[2][131] = 14'b11111111111111;
	assign font[3][131] = 14'b11111111111111;
	assign font[4][131] = 14'b11111111111111;
	assign font[5][131] = 14'b11111111111111;
	assign font[6][131] = 14'b11111111111111;
	assign font[7][131] = 14'b11111111111111;
	assign font[8][131] = 14'b11111111111111;
	assign font[9][131] = 14'b11111111111111;
	assign font[10][131] = 14'b11111111111111;
	assign font[11][131] = 14'b11111111111111;
	assign font[12][131] = 14'b11111111111111;
	assign font[13][131] = 14'b11111111111111;
	assign font[14][131] = 14'b11111111111111;
	assign font[15][131] = 14'b11111111111111;
	assign font[16][131] = 14'b11111111111111;
	assign font[17][131] = 14'b11111111111111;
	assign font[18][131] = 14'b11111111111111;
	assign font[19][131] = 14'b11111111111111;
	assign font[20][131] = 14'b11111111111111;
	assign font[21][131] = 14'b11111111111111;
	assign font[22][131] = 14'b11111111111111;
	assign font[23][131] = 14'b11111111111111;
	assign font[24][131] = 14'b11111111111111;
	assign font[25][131] = 14'b11111111111111;
	assign font[26][131] = 14'b11111111111111;
	assign font[27][131] = 14'b11111111111111;
	assign font[28][131] = 14'b11111111111111;
	assign font[29][131] = 14'b11111111111111;
	assign font[30][131] = 14'b11111111111111;
	assign font[31][131] = 14'b11111111111111;

	assign font[0][132] = 14'b11111111111111;
	assign font[1][132] = 14'b11111111111111;
	assign font[2][132] = 14'b11111111111111;
	assign font[3][132] = 14'b11111111111111;
	assign font[4][132] = 14'b11111111111111;
	assign font[5][132] = 14'b11111111111111;
	assign font[6][132] = 14'b11111111111111;
	assign font[7][132] = 14'b11111111111111;
	assign font[8][132] = 14'b11111111111111;
	assign font[9][132] = 14'b11111111111111;
	assign font[10][132] = 14'b11111111111111;
	assign font[11][132] = 14'b11111111111111;
	assign font[12][132] = 14'b11111111111111;
	assign font[13][132] = 14'b11111111111111;
	assign font[14][132] = 14'b11111111111111;
	assign font[15][132] = 14'b11111111111111;
	assign font[16][132] = 14'b11111111111111;
	assign font[17][132] = 14'b11111111111111;
	assign font[18][132] = 14'b11111111111111;
	assign font[19][132] = 14'b11111111111111;
	assign font[20][132] = 14'b11111111111111;
	assign font[21][132] = 14'b11111111111111;
	assign font[22][132] = 14'b11111111111111;
	assign font[23][132] = 14'b11111111111111;
	assign font[24][132] = 14'b11111111111111;
	assign font[25][132] = 14'b11111111111111;
	assign font[26][132] = 14'b11111111111111;
	assign font[27][132] = 14'b11111111111111;
	assign font[28][132] = 14'b11111111111111;
	assign font[29][132] = 14'b11111111111111;
	assign font[30][132] = 14'b11111111111111;
	assign font[31][132] = 14'b11111111111111;

	assign font[0][133] = 14'b11111111111111;
	assign font[1][133] = 14'b11111111111111;
	assign font[2][133] = 14'b11111111111111;
	assign font[3][133] = 14'b11111111111111;
	assign font[4][133] = 14'b11111111111111;
	assign font[5][133] = 14'b11111111111111;
	assign font[6][133] = 14'b11111111111111;
	assign font[7][133] = 14'b11111111111111;
	assign font[8][133] = 14'b11111111111111;
	assign font[9][133] = 14'b11111111111111;
	assign font[10][133] = 14'b11111111111111;
	assign font[11][133] = 14'b11111111111111;
	assign font[12][133] = 14'b11111111111111;
	assign font[13][133] = 14'b11111111111111;
	assign font[14][133] = 14'b11111111111111;
	assign font[15][133] = 14'b11111111111111;
	assign font[16][133] = 14'b11111111111111;
	assign font[17][133] = 14'b11111111111111;
	assign font[18][133] = 14'b11111111111111;
	assign font[19][133] = 14'b11111111111111;
	assign font[20][133] = 14'b11111111111111;
	assign font[21][133] = 14'b11111111111111;
	assign font[22][133] = 14'b11111111111111;
	assign font[23][133] = 14'b11111111111111;
	assign font[24][133] = 14'b11111111111111;
	assign font[25][133] = 14'b11111111111111;
	assign font[26][133] = 14'b11111111111111;
	assign font[27][133] = 14'b11111111111111;
	assign font[28][133] = 14'b11111111111111;
	assign font[29][133] = 14'b11111111111111;
	assign font[30][133] = 14'b11111111111111;
	assign font[31][133] = 14'b11111111111111;

	assign font[0][134] = 14'b11111111111111;
	assign font[1][134] = 14'b11111111111111;
	assign font[2][134] = 14'b11111111111111;
	assign font[3][134] = 14'b11111111111111;
	assign font[4][134] = 14'b11111111111111;
	assign font[5][134] = 14'b11111111111111;
	assign font[6][134] = 14'b11111111111111;
	assign font[7][134] = 14'b11111111111111;
	assign font[8][134] = 14'b11111111111111;
	assign font[9][134] = 14'b11111111111111;
	assign font[10][134] = 14'b11111111111111;
	assign font[11][134] = 14'b11111111111111;
	assign font[12][134] = 14'b11111111111111;
	assign font[13][134] = 14'b11111111111111;
	assign font[14][134] = 14'b11111111111111;
	assign font[15][134] = 14'b11111111111111;
	assign font[16][134] = 14'b11111111111111;
	assign font[17][134] = 14'b11111111111111;
	assign font[18][134] = 14'b11111111111111;
	assign font[19][134] = 14'b11111111111111;
	assign font[20][134] = 14'b11111111111111;
	assign font[21][134] = 14'b11111111111111;
	assign font[22][134] = 14'b11111111111111;
	assign font[23][134] = 14'b11111111111111;
	assign font[24][134] = 14'b11111111111111;
	assign font[25][134] = 14'b11111111111111;
	assign font[26][134] = 14'b11111111111111;
	assign font[27][134] = 14'b11111111111111;
	assign font[28][134] = 14'b11111111111111;
	assign font[29][134] = 14'b11111111111111;
	assign font[30][134] = 14'b11111111111111;
	assign font[31][134] = 14'b11111111111111;

	assign font[0][135] = 14'b11111111111111;
	assign font[1][135] = 14'b11111111111111;
	assign font[2][135] = 14'b11111111111111;
	assign font[3][135] = 14'b11111111111111;
	assign font[4][135] = 14'b11111111111111;
	assign font[5][135] = 14'b11111111111111;
	assign font[6][135] = 14'b11111111111111;
	assign font[7][135] = 14'b11111111111111;
	assign font[8][135] = 14'b11111111111111;
	assign font[9][135] = 14'b11111111111111;
	assign font[10][135] = 14'b11111111111111;
	assign font[11][135] = 14'b11111111111111;
	assign font[12][135] = 14'b11111111111111;
	assign font[13][135] = 14'b11111111111111;
	assign font[14][135] = 14'b11111111111111;
	assign font[15][135] = 14'b11111111111111;
	assign font[16][135] = 14'b11111111111111;
	assign font[17][135] = 14'b11111111111111;
	assign font[18][135] = 14'b11111111111111;
	assign font[19][135] = 14'b11111111111111;
	assign font[20][135] = 14'b11111111111111;
	assign font[21][135] = 14'b11111111111111;
	assign font[22][135] = 14'b11111111111111;
	assign font[23][135] = 14'b11111111111111;
	assign font[24][135] = 14'b11111111111111;
	assign font[25][135] = 14'b11111111111111;
	assign font[26][135] = 14'b11111111111111;
	assign font[27][135] = 14'b11111111111111;
	assign font[28][135] = 14'b11111111111111;
	assign font[29][135] = 14'b11111111111111;
	assign font[30][135] = 14'b11111111111111;
	assign font[31][135] = 14'b11111111111111;

	assign font[0][136] = 14'b11111111111111;
	assign font[1][136] = 14'b11111111111111;
	assign font[2][136] = 14'b11111111111111;
	assign font[3][136] = 14'b11111111111111;
	assign font[4][136] = 14'b11111111111111;
	assign font[5][136] = 14'b11111111111111;
	assign font[6][136] = 14'b11111111111111;
	assign font[7][136] = 14'b11111111111111;
	assign font[8][136] = 14'b11111111111111;
	assign font[9][136] = 14'b11111111111111;
	assign font[10][136] = 14'b11111111111111;
	assign font[11][136] = 14'b11111111111111;
	assign font[12][136] = 14'b11111111111111;
	assign font[13][136] = 14'b11111111111111;
	assign font[14][136] = 14'b11111111111111;
	assign font[15][136] = 14'b11111111111111;
	assign font[16][136] = 14'b11111111111111;
	assign font[17][136] = 14'b11111111111111;
	assign font[18][136] = 14'b11111111111111;
	assign font[19][136] = 14'b11111111111111;
	assign font[20][136] = 14'b11111111111111;
	assign font[21][136] = 14'b11111111111111;
	assign font[22][136] = 14'b11111111111111;
	assign font[23][136] = 14'b11111111111111;
	assign font[24][136] = 14'b11111111111111;
	assign font[25][136] = 14'b11111111111111;
	assign font[26][136] = 14'b11111111111111;
	assign font[27][136] = 14'b11111111111111;
	assign font[28][136] = 14'b11111111111111;
	assign font[29][136] = 14'b11111111111111;
	assign font[30][136] = 14'b11111111111111;
	assign font[31][136] = 14'b11111111111111;

	assign font[0][137] = 14'b11111111111111;
	assign font[1][137] = 14'b11111111111111;
	assign font[2][137] = 14'b11111111111111;
	assign font[3][137] = 14'b11111111111111;
	assign font[4][137] = 14'b11111111111111;
	assign font[5][137] = 14'b11111111111111;
	assign font[6][137] = 14'b11111111111111;
	assign font[7][137] = 14'b11111111111111;
	assign font[8][137] = 14'b11111111111111;
	assign font[9][137] = 14'b11111111111111;
	assign font[10][137] = 14'b11111111111111;
	assign font[11][137] = 14'b11111111111111;
	assign font[12][137] = 14'b11111111111111;
	assign font[13][137] = 14'b11111111111111;
	assign font[14][137] = 14'b11111111111111;
	assign font[15][137] = 14'b11111111111111;
	assign font[16][137] = 14'b11111111111111;
	assign font[17][137] = 14'b11111111111111;
	assign font[18][137] = 14'b11111111111111;
	assign font[19][137] = 14'b11111111111111;
	assign font[20][137] = 14'b11111111111111;
	assign font[21][137] = 14'b11111111111111;
	assign font[22][137] = 14'b11111111111111;
	assign font[23][137] = 14'b11111111111111;
	assign font[24][137] = 14'b11111111111111;
	assign font[25][137] = 14'b11111111111111;
	assign font[26][137] = 14'b11111111111111;
	assign font[27][137] = 14'b11111111111111;
	assign font[28][137] = 14'b11111111111111;
	assign font[29][137] = 14'b11111111111111;
	assign font[30][137] = 14'b11111111111111;
	assign font[31][137] = 14'b11111111111111;

	assign font[0][138] = 14'b11111111111111;
	assign font[1][138] = 14'b11111111111111;
	assign font[2][138] = 14'b11111111111111;
	assign font[3][138] = 14'b11111111111111;
	assign font[4][138] = 14'b11111111111111;
	assign font[5][138] = 14'b11111111111111;
	assign font[6][138] = 14'b11111111111111;
	assign font[7][138] = 14'b11111111111111;
	assign font[8][138] = 14'b11111111111111;
	assign font[9][138] = 14'b11111111111111;
	assign font[10][138] = 14'b11111111111111;
	assign font[11][138] = 14'b11111111111111;
	assign font[12][138] = 14'b11111111111111;
	assign font[13][138] = 14'b11111111111111;
	assign font[14][138] = 14'b11111111111111;
	assign font[15][138] = 14'b11111111111111;
	assign font[16][138] = 14'b11111111111111;
	assign font[17][138] = 14'b11111111111111;
	assign font[18][138] = 14'b11111111111111;
	assign font[19][138] = 14'b11111111111111;
	assign font[20][138] = 14'b11111111111111;
	assign font[21][138] = 14'b11111111111111;
	assign font[22][138] = 14'b11111111111111;
	assign font[23][138] = 14'b11111111111111;
	assign font[24][138] = 14'b11111111111111;
	assign font[25][138] = 14'b11111111111111;
	assign font[26][138] = 14'b11111111111111;
	assign font[27][138] = 14'b11111111111111;
	assign font[28][138] = 14'b11111111111111;
	assign font[29][138] = 14'b11111111111111;
	assign font[30][138] = 14'b11111111111111;
	assign font[31][138] = 14'b11111111111111;

	assign font[0][139] = 14'b11111111111111;
	assign font[1][139] = 14'b11111111111111;
	assign font[2][139] = 14'b11111111111111;
	assign font[3][139] = 14'b11111111111111;
	assign font[4][139] = 14'b11111111111111;
	assign font[5][139] = 14'b11111111111111;
	assign font[6][139] = 14'b11111111111111;
	assign font[7][139] = 14'b11111111111111;
	assign font[8][139] = 14'b11111111111111;
	assign font[9][139] = 14'b11111111111111;
	assign font[10][139] = 14'b11111111111111;
	assign font[11][139] = 14'b11111111111111;
	assign font[12][139] = 14'b11111111111111;
	assign font[13][139] = 14'b11111111111111;
	assign font[14][139] = 14'b11111111111111;
	assign font[15][139] = 14'b11111111111111;
	assign font[16][139] = 14'b11111111111111;
	assign font[17][139] = 14'b11111111111111;
	assign font[18][139] = 14'b11111111111111;
	assign font[19][139] = 14'b11111111111111;
	assign font[20][139] = 14'b11111111111111;
	assign font[21][139] = 14'b11111111111111;
	assign font[22][139] = 14'b11111111111111;
	assign font[23][139] = 14'b11111111111111;
	assign font[24][139] = 14'b11111111111111;
	assign font[25][139] = 14'b11111111111111;
	assign font[26][139] = 14'b11111111111111;
	assign font[27][139] = 14'b11111111111111;
	assign font[28][139] = 14'b11111111111111;
	assign font[29][139] = 14'b11111111111111;
	assign font[30][139] = 14'b11111111111111;
	assign font[31][139] = 14'b11111111111111;

	assign font[0][140] = 14'b11111111111111;
	assign font[1][140] = 14'b11111111111111;
	assign font[2][140] = 14'b11111111111111;
	assign font[3][140] = 14'b11111111111111;
	assign font[4][140] = 14'b11111111111111;
	assign font[5][140] = 14'b11111111111111;
	assign font[6][140] = 14'b11111111111111;
	assign font[7][140] = 14'b11111111111111;
	assign font[8][140] = 14'b11111111111111;
	assign font[9][140] = 14'b11111111111111;
	assign font[10][140] = 14'b11111111111111;
	assign font[11][140] = 14'b11111111111111;
	assign font[12][140] = 14'b11111111111111;
	assign font[13][140] = 14'b11111111111111;
	assign font[14][140] = 14'b11111111111111;
	assign font[15][140] = 14'b11111111111111;
	assign font[16][140] = 14'b11111111111111;
	assign font[17][140] = 14'b11111111111111;
	assign font[18][140] = 14'b11111111111111;
	assign font[19][140] = 14'b11111111111111;
	assign font[20][140] = 14'b11111111111111;
	assign font[21][140] = 14'b11111111111111;
	assign font[22][140] = 14'b11111111111111;
	assign font[23][140] = 14'b11111111111111;
	assign font[24][140] = 14'b11111111111111;
	assign font[25][140] = 14'b11111111111111;
	assign font[26][140] = 14'b11111111111111;
	assign font[27][140] = 14'b11111111111111;
	assign font[28][140] = 14'b11111111111111;
	assign font[29][140] = 14'b11111111111111;
	assign font[30][140] = 14'b11111111111111;
	assign font[31][140] = 14'b11111111111111;

	assign font[0][141] = 14'b11111111111111;
	assign font[1][141] = 14'b11111111111111;
	assign font[2][141] = 14'b11111111111111;
	assign font[3][141] = 14'b11111111111111;
	assign font[4][141] = 14'b11111111111111;
	assign font[5][141] = 14'b11111111111111;
	assign font[6][141] = 14'b11111111111111;
	assign font[7][141] = 14'b11111111111111;
	assign font[8][141] = 14'b11111111111111;
	assign font[9][141] = 14'b11111111111111;
	assign font[10][141] = 14'b11111111111111;
	assign font[11][141] = 14'b11111111111111;
	assign font[12][141] = 14'b11111111111111;
	assign font[13][141] = 14'b11111111111111;
	assign font[14][141] = 14'b11111111111111;
	assign font[15][141] = 14'b11111111111111;
	assign font[16][141] = 14'b11111111111111;
	assign font[17][141] = 14'b11111111111111;
	assign font[18][141] = 14'b11111111111111;
	assign font[19][141] = 14'b11111111111111;
	assign font[20][141] = 14'b11111111111111;
	assign font[21][141] = 14'b11111111111111;
	assign font[22][141] = 14'b11111111111111;
	assign font[23][141] = 14'b11111111111111;
	assign font[24][141] = 14'b11111111111111;
	assign font[25][141] = 14'b11111111111111;
	assign font[26][141] = 14'b11111111111111;
	assign font[27][141] = 14'b11111111111111;
	assign font[28][141] = 14'b11111111111111;
	assign font[29][141] = 14'b11111111111111;
	assign font[30][141] = 14'b11111111111111;
	assign font[31][141] = 14'b11111111111111;

	assign font[0][142] = 14'b11111111111111;
	assign font[1][142] = 14'b11111111111111;
	assign font[2][142] = 14'b11111111111111;
	assign font[3][142] = 14'b11111111111111;
	assign font[4][142] = 14'b11111111111111;
	assign font[5][142] = 14'b11111111111111;
	assign font[6][142] = 14'b11111111111111;
	assign font[7][142] = 14'b11111111111111;
	assign font[8][142] = 14'b11111111111111;
	assign font[9][142] = 14'b11111111111111;
	assign font[10][142] = 14'b11111111111111;
	assign font[11][142] = 14'b11111111111111;
	assign font[12][142] = 14'b11111111111111;
	assign font[13][142] = 14'b11111111111111;
	assign font[14][142] = 14'b11111111111111;
	assign font[15][142] = 14'b11111111111111;
	assign font[16][142] = 14'b11111111111111;
	assign font[17][142] = 14'b11111111111111;
	assign font[18][142] = 14'b11111111111111;
	assign font[19][142] = 14'b11111111111111;
	assign font[20][142] = 14'b11111111111111;
	assign font[21][142] = 14'b11111111111111;
	assign font[22][142] = 14'b11111111111111;
	assign font[23][142] = 14'b11111111111111;
	assign font[24][142] = 14'b11111111111111;
	assign font[25][142] = 14'b11111111111111;
	assign font[26][142] = 14'b11111111111111;
	assign font[27][142] = 14'b11111111111111;
	assign font[28][142] = 14'b11111111111111;
	assign font[29][142] = 14'b11111111111111;
	assign font[30][142] = 14'b11111111111111;
	assign font[31][142] = 14'b11111111111111;

	assign font[0][143] = 14'b11111111111111;
	assign font[1][143] = 14'b11111111111111;
	assign font[2][143] = 14'b11111111111111;
	assign font[3][143] = 14'b11111111111111;
	assign font[4][143] = 14'b11111111111111;
	assign font[5][143] = 14'b11111111111111;
	assign font[6][143] = 14'b11111111111111;
	assign font[7][143] = 14'b11111111111111;
	assign font[8][143] = 14'b11111111111111;
	assign font[9][143] = 14'b11111111111111;
	assign font[10][143] = 14'b11111111111111;
	assign font[11][143] = 14'b11111111111111;
	assign font[12][143] = 14'b11111111111111;
	assign font[13][143] = 14'b11111111111111;
	assign font[14][143] = 14'b11111111111111;
	assign font[15][143] = 14'b11111111111111;
	assign font[16][143] = 14'b11111111111111;
	assign font[17][143] = 14'b11111111111111;
	assign font[18][143] = 14'b11111111111111;
	assign font[19][143] = 14'b11111111111111;
	assign font[20][143] = 14'b11111111111111;
	assign font[21][143] = 14'b11111111111111;
	assign font[22][143] = 14'b11111111111111;
	assign font[23][143] = 14'b11111111111111;
	assign font[24][143] = 14'b11111111111111;
	assign font[25][143] = 14'b11111111111111;
	assign font[26][143] = 14'b11111111111111;
	assign font[27][143] = 14'b11111111111111;
	assign font[28][143] = 14'b11111111111111;
	assign font[29][143] = 14'b11111111111111;
	assign font[30][143] = 14'b11111111111111;
	assign font[31][143] = 14'b11111111111111;

	assign font[0][144] = 14'b11111111111111;
	assign font[1][144] = 14'b11111111111111;
	assign font[2][144] = 14'b11111111111111;
	assign font[3][144] = 14'b11111111111111;
	assign font[4][144] = 14'b11111111111111;
	assign font[5][144] = 14'b11111111111111;
	assign font[6][144] = 14'b11111111111111;
	assign font[7][144] = 14'b11111111111111;
	assign font[8][144] = 14'b11111111111111;
	assign font[9][144] = 14'b11111111111111;
	assign font[10][144] = 14'b11111111111111;
	assign font[11][144] = 14'b11111111111111;
	assign font[12][144] = 14'b11111111111111;
	assign font[13][144] = 14'b11111111111111;
	assign font[14][144] = 14'b11111111111111;
	assign font[15][144] = 14'b11111111111111;
	assign font[16][144] = 14'b11111111111111;
	assign font[17][144] = 14'b11111111111111;
	assign font[18][144] = 14'b11111111111111;
	assign font[19][144] = 14'b11111111111111;
	assign font[20][144] = 14'b11111111111111;
	assign font[21][144] = 14'b11111111111111;
	assign font[22][144] = 14'b11111111111111;
	assign font[23][144] = 14'b11111111111111;
	assign font[24][144] = 14'b11111111111111;
	assign font[25][144] = 14'b11111111111111;
	assign font[26][144] = 14'b11111111111111;
	assign font[27][144] = 14'b11111111111111;
	assign font[28][144] = 14'b11111111111111;
	assign font[29][144] = 14'b11111111111111;
	assign font[30][144] = 14'b11111111111111;
	assign font[31][144] = 14'b11111111111111;

	assign font[0][145] = 14'b11111111111111;
	assign font[1][145] = 14'b11111111111111;
	assign font[2][145] = 14'b11111111111111;
	assign font[3][145] = 14'b11111111111111;
	assign font[4][145] = 14'b11111111111111;
	assign font[5][145] = 14'b11111111111111;
	assign font[6][145] = 14'b11111111111111;
	assign font[7][145] = 14'b11111111111111;
	assign font[8][145] = 14'b11111111111111;
	assign font[9][145] = 14'b11111111111111;
	assign font[10][145] = 14'b11111111111111;
	assign font[11][145] = 14'b11111111111111;
	assign font[12][145] = 14'b11111111111111;
	assign font[13][145] = 14'b11111111111111;
	assign font[14][145] = 14'b11111111111111;
	assign font[15][145] = 14'b11111111111111;
	assign font[16][145] = 14'b11111111111111;
	assign font[17][145] = 14'b11111111111111;
	assign font[18][145] = 14'b11111111111111;
	assign font[19][145] = 14'b11111111111111;
	assign font[20][145] = 14'b11111111111111;
	assign font[21][145] = 14'b11111111111111;
	assign font[22][145] = 14'b11111111111111;
	assign font[23][145] = 14'b11111111111111;
	assign font[24][145] = 14'b11111111111111;
	assign font[25][145] = 14'b11111111111111;
	assign font[26][145] = 14'b11111111111111;
	assign font[27][145] = 14'b11111111111111;
	assign font[28][145] = 14'b11111111111111;
	assign font[29][145] = 14'b11111111111111;
	assign font[30][145] = 14'b11111111111111;
	assign font[31][145] = 14'b11111111111111;

	assign font[0][146] = 14'b11111111111111;
	assign font[1][146] = 14'b11111111111111;
	assign font[2][146] = 14'b11111111111111;
	assign font[3][146] = 14'b11111111111111;
	assign font[4][146] = 14'b11111111111111;
	assign font[5][146] = 14'b11111111111111;
	assign font[6][146] = 14'b11111111111111;
	assign font[7][146] = 14'b11111111111111;
	assign font[8][146] = 14'b11111111111111;
	assign font[9][146] = 14'b11111111111111;
	assign font[10][146] = 14'b11111111111111;
	assign font[11][146] = 14'b11111111111111;
	assign font[12][146] = 14'b11111111111111;
	assign font[13][146] = 14'b11111111111111;
	assign font[14][146] = 14'b11111111111111;
	assign font[15][146] = 14'b11111111111111;
	assign font[16][146] = 14'b11111111111111;
	assign font[17][146] = 14'b11111111111111;
	assign font[18][146] = 14'b11111111111111;
	assign font[19][146] = 14'b11111111111111;
	assign font[20][146] = 14'b11111111111111;
	assign font[21][146] = 14'b11111111111111;
	assign font[22][146] = 14'b11111111111111;
	assign font[23][146] = 14'b11111111111111;
	assign font[24][146] = 14'b11111111111111;
	assign font[25][146] = 14'b11111111111111;
	assign font[26][146] = 14'b11111111111111;
	assign font[27][146] = 14'b11111111111111;
	assign font[28][146] = 14'b11111111111111;
	assign font[29][146] = 14'b11111111111111;
	assign font[30][146] = 14'b11111111111111;
	assign font[31][146] = 14'b11111111111111;

	assign font[0][147] = 14'b11111111111111;
	assign font[1][147] = 14'b11111111111111;
	assign font[2][147] = 14'b11111111111111;
	assign font[3][147] = 14'b11111111111111;
	assign font[4][147] = 14'b11111111111111;
	assign font[5][147] = 14'b11111111111111;
	assign font[6][147] = 14'b11111111111111;
	assign font[7][147] = 14'b11111111111111;
	assign font[8][147] = 14'b11111111111111;
	assign font[9][147] = 14'b11111111111111;
	assign font[10][147] = 14'b11111111111111;
	assign font[11][147] = 14'b11111111111111;
	assign font[12][147] = 14'b11111111111111;
	assign font[13][147] = 14'b11111111111111;
	assign font[14][147] = 14'b11111111111111;
	assign font[15][147] = 14'b11111111111111;
	assign font[16][147] = 14'b11111111111111;
	assign font[17][147] = 14'b11111111111111;
	assign font[18][147] = 14'b11111111111111;
	assign font[19][147] = 14'b11111111111111;
	assign font[20][147] = 14'b11111111111111;
	assign font[21][147] = 14'b11111111111111;
	assign font[22][147] = 14'b11111111111111;
	assign font[23][147] = 14'b11111111111111;
	assign font[24][147] = 14'b11111111111111;
	assign font[25][147] = 14'b11111111111111;
	assign font[26][147] = 14'b11111111111111;
	assign font[27][147] = 14'b11111111111111;
	assign font[28][147] = 14'b11111111111111;
	assign font[29][147] = 14'b11111111111111;
	assign font[30][147] = 14'b11111111111111;
	assign font[31][147] = 14'b11111111111111;

	assign font[0][148] = 14'b11111111111111;
	assign font[1][148] = 14'b11111111111111;
	assign font[2][148] = 14'b11111111111111;
	assign font[3][148] = 14'b11111111111111;
	assign font[4][148] = 14'b11111111111111;
	assign font[5][148] = 14'b11111111111111;
	assign font[6][148] = 14'b11111111111111;
	assign font[7][148] = 14'b11111111111111;
	assign font[8][148] = 14'b11111111111111;
	assign font[9][148] = 14'b11111111111111;
	assign font[10][148] = 14'b11111111111111;
	assign font[11][148] = 14'b11111111111111;
	assign font[12][148] = 14'b11111111111111;
	assign font[13][148] = 14'b11111111111111;
	assign font[14][148] = 14'b11111111111111;
	assign font[15][148] = 14'b11111111111111;
	assign font[16][148] = 14'b11111111111111;
	assign font[17][148] = 14'b11111111111111;
	assign font[18][148] = 14'b11111111111111;
	assign font[19][148] = 14'b11111111111111;
	assign font[20][148] = 14'b11111111111111;
	assign font[21][148] = 14'b11111111111111;
	assign font[22][148] = 14'b11111111111111;
	assign font[23][148] = 14'b11111111111111;
	assign font[24][148] = 14'b11111111111111;
	assign font[25][148] = 14'b11111111111111;
	assign font[26][148] = 14'b11111111111111;
	assign font[27][148] = 14'b11111111111111;
	assign font[28][148] = 14'b11111111111111;
	assign font[29][148] = 14'b11111111111111;
	assign font[30][148] = 14'b11111111111111;
	assign font[31][148] = 14'b11111111111111;

	assign font[0][149] = 14'b11111111111111;
	assign font[1][149] = 14'b11111111111111;
	assign font[2][149] = 14'b11111111111111;
	assign font[3][149] = 14'b11111111111111;
	assign font[4][149] = 14'b11111111111111;
	assign font[5][149] = 14'b11111111111111;
	assign font[6][149] = 14'b11111111111111;
	assign font[7][149] = 14'b11111111111111;
	assign font[8][149] = 14'b11111111111111;
	assign font[9][149] = 14'b11111111111111;
	assign font[10][149] = 14'b11111111111111;
	assign font[11][149] = 14'b11111111111111;
	assign font[12][149] = 14'b11111111111111;
	assign font[13][149] = 14'b11111111111111;
	assign font[14][149] = 14'b11111111111111;
	assign font[15][149] = 14'b11111111111111;
	assign font[16][149] = 14'b11111111111111;
	assign font[17][149] = 14'b11111111111111;
	assign font[18][149] = 14'b11111111111111;
	assign font[19][149] = 14'b11111111111111;
	assign font[20][149] = 14'b11111111111111;
	assign font[21][149] = 14'b11111111111111;
	assign font[22][149] = 14'b11111111111111;
	assign font[23][149] = 14'b11111111111111;
	assign font[24][149] = 14'b11111111111111;
	assign font[25][149] = 14'b11111111111111;
	assign font[26][149] = 14'b11111111111111;
	assign font[27][149] = 14'b11111111111111;
	assign font[28][149] = 14'b11111111111111;
	assign font[29][149] = 14'b11111111111111;
	assign font[30][149] = 14'b11111111111111;
	assign font[31][149] = 14'b11111111111111;

	assign font[0][150] = 14'b11111111111111;
	assign font[1][150] = 14'b11111111111111;
	assign font[2][150] = 14'b11111111111111;
	assign font[3][150] = 14'b11111111111111;
	assign font[4][150] = 14'b11111111111111;
	assign font[5][150] = 14'b11111111111111;
	assign font[6][150] = 14'b11111111111111;
	assign font[7][150] = 14'b11111111111111;
	assign font[8][150] = 14'b11111111111111;
	assign font[9][150] = 14'b11111111111111;
	assign font[10][150] = 14'b11111111111111;
	assign font[11][150] = 14'b11111111111111;
	assign font[12][150] = 14'b11111111111111;
	assign font[13][150] = 14'b11111111111111;
	assign font[14][150] = 14'b11111111111111;
	assign font[15][150] = 14'b11111111111111;
	assign font[16][150] = 14'b11111111111111;
	assign font[17][150] = 14'b11111111111111;
	assign font[18][150] = 14'b11111111111111;
	assign font[19][150] = 14'b11111111111111;
	assign font[20][150] = 14'b11111111111111;
	assign font[21][150] = 14'b11111111111111;
	assign font[22][150] = 14'b11111111111111;
	assign font[23][150] = 14'b11111111111111;
	assign font[24][150] = 14'b11111111111111;
	assign font[25][150] = 14'b11111111111111;
	assign font[26][150] = 14'b11111111111111;
	assign font[27][150] = 14'b11111111111111;
	assign font[28][150] = 14'b11111111111111;
	assign font[29][150] = 14'b11111111111111;
	assign font[30][150] = 14'b11111111111111;
	assign font[31][150] = 14'b11111111111111;

	assign font[0][151] = 14'b11111111111111;
	assign font[1][151] = 14'b11111111111111;
	assign font[2][151] = 14'b11111111111111;
	assign font[3][151] = 14'b11111111111111;
	assign font[4][151] = 14'b11111111111111;
	assign font[5][151] = 14'b11111111111111;
	assign font[6][151] = 14'b11111111111111;
	assign font[7][151] = 14'b11111111111111;
	assign font[8][151] = 14'b11111111111111;
	assign font[9][151] = 14'b11111111111111;
	assign font[10][151] = 14'b11111111111111;
	assign font[11][151] = 14'b11111111111111;
	assign font[12][151] = 14'b11111111111111;
	assign font[13][151] = 14'b11111111111111;
	assign font[14][151] = 14'b11111111111111;
	assign font[15][151] = 14'b11111111111111;
	assign font[16][151] = 14'b11111111111111;
	assign font[17][151] = 14'b11111111111111;
	assign font[18][151] = 14'b11111111111111;
	assign font[19][151] = 14'b11111111111111;
	assign font[20][151] = 14'b11111111111111;
	assign font[21][151] = 14'b11111111111111;
	assign font[22][151] = 14'b11111111111111;
	assign font[23][151] = 14'b11111111111111;
	assign font[24][151] = 14'b11111111111111;
	assign font[25][151] = 14'b11111111111111;
	assign font[26][151] = 14'b11111111111111;
	assign font[27][151] = 14'b11111111111111;
	assign font[28][151] = 14'b11111111111111;
	assign font[29][151] = 14'b11111111111111;
	assign font[30][151] = 14'b11111111111111;
	assign font[31][151] = 14'b11111111111111;

	assign font[0][152] = 14'b11111111111111;
	assign font[1][152] = 14'b11111111111111;
	assign font[2][152] = 14'b11111111111111;
	assign font[3][152] = 14'b11111111111111;
	assign font[4][152] = 14'b11111111111111;
	assign font[5][152] = 14'b11111111111111;
	assign font[6][152] = 14'b11111111111111;
	assign font[7][152] = 14'b11111111111111;
	assign font[8][152] = 14'b11111111111111;
	assign font[9][152] = 14'b11111111111111;
	assign font[10][152] = 14'b11111111111111;
	assign font[11][152] = 14'b11111111111111;
	assign font[12][152] = 14'b11111111111111;
	assign font[13][152] = 14'b11111111111111;
	assign font[14][152] = 14'b11111111111111;
	assign font[15][152] = 14'b11111111111111;
	assign font[16][152] = 14'b11111111111111;
	assign font[17][152] = 14'b11111111111111;
	assign font[18][152] = 14'b11111111111111;
	assign font[19][152] = 14'b11111111111111;
	assign font[20][152] = 14'b11111111111111;
	assign font[21][152] = 14'b11111111111111;
	assign font[22][152] = 14'b11111111111111;
	assign font[23][152] = 14'b11111111111111;
	assign font[24][152] = 14'b11111111111111;
	assign font[25][152] = 14'b11111111111111;
	assign font[26][152] = 14'b11111111111111;
	assign font[27][152] = 14'b11111111111111;
	assign font[28][152] = 14'b11111111111111;
	assign font[29][152] = 14'b11111111111111;
	assign font[30][152] = 14'b11111111111111;
	assign font[31][152] = 14'b11111111111111;

	assign font[0][153] = 14'b11111111111111;
	assign font[1][153] = 14'b11111111111111;
	assign font[2][153] = 14'b11111111111111;
	assign font[3][153] = 14'b11111111111111;
	assign font[4][153] = 14'b11111111111111;
	assign font[5][153] = 14'b11111111111111;
	assign font[6][153] = 14'b11111111111111;
	assign font[7][153] = 14'b11111111111111;
	assign font[8][153] = 14'b11111111111111;
	assign font[9][153] = 14'b11111111111111;
	assign font[10][153] = 14'b11111111111111;
	assign font[11][153] = 14'b11111111111111;
	assign font[12][153] = 14'b11111111111111;
	assign font[13][153] = 14'b11111111111111;
	assign font[14][153] = 14'b11111111111111;
	assign font[15][153] = 14'b11111111111111;
	assign font[16][153] = 14'b11111111111111;
	assign font[17][153] = 14'b11111111111111;
	assign font[18][153] = 14'b11111111111111;
	assign font[19][153] = 14'b11111111111111;
	assign font[20][153] = 14'b11111111111111;
	assign font[21][153] = 14'b11111111111111;
	assign font[22][153] = 14'b11111111111111;
	assign font[23][153] = 14'b11111111111111;
	assign font[24][153] = 14'b11111111111111;
	assign font[25][153] = 14'b11111111111111;
	assign font[26][153] = 14'b11111111111111;
	assign font[27][153] = 14'b11111111111111;
	assign font[28][153] = 14'b11111111111111;
	assign font[29][153] = 14'b11111111111111;
	assign font[30][153] = 14'b11111111111111;
	assign font[31][153] = 14'b11111111111111;

	assign font[0][154] = 14'b11111111111111;
	assign font[1][154] = 14'b11111111111111;
	assign font[2][154] = 14'b11111111111111;
	assign font[3][154] = 14'b11111111111111;
	assign font[4][154] = 14'b11111111111111;
	assign font[5][154] = 14'b11111111111111;
	assign font[6][154] = 14'b11111111111111;
	assign font[7][154] = 14'b11111111111111;
	assign font[8][154] = 14'b11111111111111;
	assign font[9][154] = 14'b11111111111111;
	assign font[10][154] = 14'b11111111111111;
	assign font[11][154] = 14'b11111111111111;
	assign font[12][154] = 14'b11111111111111;
	assign font[13][154] = 14'b11111111111111;
	assign font[14][154] = 14'b11111111111111;
	assign font[15][154] = 14'b11111111111111;
	assign font[16][154] = 14'b11111111111111;
	assign font[17][154] = 14'b11111111111111;
	assign font[18][154] = 14'b11111111111111;
	assign font[19][154] = 14'b11111111111111;
	assign font[20][154] = 14'b11111111111111;
	assign font[21][154] = 14'b11111111111111;
	assign font[22][154] = 14'b11111111111111;
	assign font[23][154] = 14'b11111111111111;
	assign font[24][154] = 14'b11111111111111;
	assign font[25][154] = 14'b11111111111111;
	assign font[26][154] = 14'b11111111111111;
	assign font[27][154] = 14'b11111111111111;
	assign font[28][154] = 14'b11111111111111;
	assign font[29][154] = 14'b11111111111111;
	assign font[30][154] = 14'b11111111111111;
	assign font[31][154] = 14'b11111111111111;

	assign font[0][155] = 14'b11111111111111;
	assign font[1][155] = 14'b11111111111111;
	assign font[2][155] = 14'b11111111111111;
	assign font[3][155] = 14'b11111111111111;
	assign font[4][155] = 14'b11111111111111;
	assign font[5][155] = 14'b11111111111111;
	assign font[6][155] = 14'b11111111111111;
	assign font[7][155] = 14'b11111111111111;
	assign font[8][155] = 14'b11111111111111;
	assign font[9][155] = 14'b11111111111111;
	assign font[10][155] = 14'b11111111111111;
	assign font[11][155] = 14'b11111111111111;
	assign font[12][155] = 14'b11111111111111;
	assign font[13][155] = 14'b11111111111111;
	assign font[14][155] = 14'b11111111111111;
	assign font[15][155] = 14'b11111111111111;
	assign font[16][155] = 14'b11111111111111;
	assign font[17][155] = 14'b11111111111111;
	assign font[18][155] = 14'b11111111111111;
	assign font[19][155] = 14'b11111111111111;
	assign font[20][155] = 14'b11111111111111;
	assign font[21][155] = 14'b11111111111111;
	assign font[22][155] = 14'b11111111111111;
	assign font[23][155] = 14'b11111111111111;
	assign font[24][155] = 14'b11111111111111;
	assign font[25][155] = 14'b11111111111111;
	assign font[26][155] = 14'b11111111111111;
	assign font[27][155] = 14'b11111111111111;
	assign font[28][155] = 14'b11111111111111;
	assign font[29][155] = 14'b11111111111111;
	assign font[30][155] = 14'b11111111111111;
	assign font[31][155] = 14'b11111111111111;

	assign font[0][156] = 14'b11111111111111;
	assign font[1][156] = 14'b11111111111111;
	assign font[2][156] = 14'b11111111111111;
	assign font[3][156] = 14'b11111111111111;
	assign font[4][156] = 14'b11111111111111;
	assign font[5][156] = 14'b11111111111111;
	assign font[6][156] = 14'b11111111111111;
	assign font[7][156] = 14'b11111111111111;
	assign font[8][156] = 14'b11111111111111;
	assign font[9][156] = 14'b11111111111111;
	assign font[10][156] = 14'b11111111111111;
	assign font[11][156] = 14'b11111111111111;
	assign font[12][156] = 14'b11111111111111;
	assign font[13][156] = 14'b11111111111111;
	assign font[14][156] = 14'b11111111111111;
	assign font[15][156] = 14'b11111111111111;
	assign font[16][156] = 14'b11111111111111;
	assign font[17][156] = 14'b11111111111111;
	assign font[18][156] = 14'b11111111111111;
	assign font[19][156] = 14'b11111111111111;
	assign font[20][156] = 14'b11111111111111;
	assign font[21][156] = 14'b11111111111111;
	assign font[22][156] = 14'b11111111111111;
	assign font[23][156] = 14'b11111111111111;
	assign font[24][156] = 14'b11111111111111;
	assign font[25][156] = 14'b11111111111111;
	assign font[26][156] = 14'b11111111111111;
	assign font[27][156] = 14'b11111111111111;
	assign font[28][156] = 14'b11111111111111;
	assign font[29][156] = 14'b11111111111111;
	assign font[30][156] = 14'b11111111111111;
	assign font[31][156] = 14'b11111111111111;

	assign font[0][157] = 14'b11111111111111;
	assign font[1][157] = 14'b11111111111111;
	assign font[2][157] = 14'b11111111111111;
	assign font[3][157] = 14'b11111111111111;
	assign font[4][157] = 14'b11111111111111;
	assign font[5][157] = 14'b11111111111111;
	assign font[6][157] = 14'b11111111111111;
	assign font[7][157] = 14'b11111111111111;
	assign font[8][157] = 14'b11111111111111;
	assign font[9][157] = 14'b11111111111111;
	assign font[10][157] = 14'b11111111111111;
	assign font[11][157] = 14'b11111111111111;
	assign font[12][157] = 14'b11111111111111;
	assign font[13][157] = 14'b11111111111111;
	assign font[14][157] = 14'b11111111111111;
	assign font[15][157] = 14'b11111111111111;
	assign font[16][157] = 14'b11111111111111;
	assign font[17][157] = 14'b11111111111111;
	assign font[18][157] = 14'b11111111111111;
	assign font[19][157] = 14'b11111111111111;
	assign font[20][157] = 14'b11111111111111;
	assign font[21][157] = 14'b11111111111111;
	assign font[22][157] = 14'b11111111111111;
	assign font[23][157] = 14'b11111111111111;
	assign font[24][157] = 14'b11111111111111;
	assign font[25][157] = 14'b11111111111111;
	assign font[26][157] = 14'b11111111111111;
	assign font[27][157] = 14'b11111111111111;
	assign font[28][157] = 14'b11111111111111;
	assign font[29][157] = 14'b11111111111111;
	assign font[30][157] = 14'b11111111111111;
	assign font[31][157] = 14'b11111111111111;

	assign font[0][158] = 14'b11111111111111;
	assign font[1][158] = 14'b11111111111111;
	assign font[2][158] = 14'b11111111111111;
	assign font[3][158] = 14'b11111111111111;
	assign font[4][158] = 14'b11111111111111;
	assign font[5][158] = 14'b11111111111111;
	assign font[6][158] = 14'b11111111111111;
	assign font[7][158] = 14'b11111111111111;
	assign font[8][158] = 14'b11111111111111;
	assign font[9][158] = 14'b11111111111111;
	assign font[10][158] = 14'b11111111111111;
	assign font[11][158] = 14'b11111111111111;
	assign font[12][158] = 14'b11111111111111;
	assign font[13][158] = 14'b11111111111111;
	assign font[14][158] = 14'b11111111111111;
	assign font[15][158] = 14'b11111111111111;
	assign font[16][158] = 14'b11111111111111;
	assign font[17][158] = 14'b11111111111111;
	assign font[18][158] = 14'b11111111111111;
	assign font[19][158] = 14'b11111111111111;
	assign font[20][158] = 14'b11111111111111;
	assign font[21][158] = 14'b11111111111111;
	assign font[22][158] = 14'b11111111111111;
	assign font[23][158] = 14'b11111111111111;
	assign font[24][158] = 14'b11111111111111;
	assign font[25][158] = 14'b11111111111111;
	assign font[26][158] = 14'b11111111111111;
	assign font[27][158] = 14'b11111111111111;
	assign font[28][158] = 14'b11111111111111;
	assign font[29][158] = 14'b11111111111111;
	assign font[30][158] = 14'b11111111111111;
	assign font[31][158] = 14'b11111111111111;

	assign font[0][159] = 14'b11111111111111;
	assign font[1][159] = 14'b11111111111111;
	assign font[2][159] = 14'b11111111111111;
	assign font[3][159] = 14'b11111111111111;
	assign font[4][159] = 14'b11111111111111;
	assign font[5][159] = 14'b11111111111111;
	assign font[6][159] = 14'b11111111111111;
	assign font[7][159] = 14'b11111111111111;
	assign font[8][159] = 14'b11111111111111;
	assign font[9][159] = 14'b11111111111111;
	assign font[10][159] = 14'b11111111111111;
	assign font[11][159] = 14'b11111111111111;
	assign font[12][159] = 14'b11111111111111;
	assign font[13][159] = 14'b11111111111111;
	assign font[14][159] = 14'b11111111111111;
	assign font[15][159] = 14'b11111111111111;
	assign font[16][159] = 14'b11111111111111;
	assign font[17][159] = 14'b11111111111111;
	assign font[18][159] = 14'b11111111111111;
	assign font[19][159] = 14'b11111111111111;
	assign font[20][159] = 14'b11111111111111;
	assign font[21][159] = 14'b11111111111111;
	assign font[22][159] = 14'b11111111111111;
	assign font[23][159] = 14'b11111111111111;
	assign font[24][159] = 14'b11111111111111;
	assign font[25][159] = 14'b11111111111111;
	assign font[26][159] = 14'b11111111111111;
	assign font[27][159] = 14'b11111111111111;
	assign font[28][159] = 14'b11111111111111;
	assign font[29][159] = 14'b11111111111111;
	assign font[30][159] = 14'b11111111111111;
	assign font[31][159] = 14'b11111111111111;

	assign font[0][160] = 14'b11111111111111;
	assign font[1][160] = 14'b11111111111111;
	assign font[2][160] = 14'b11111111111111;
	assign font[3][160] = 14'b11111111111111;
	assign font[4][160] = 14'b11111111111111;
	assign font[5][160] = 14'b11111111111111;
	assign font[6][160] = 14'b11111111111111;
	assign font[7][160] = 14'b11111111111111;
	assign font[8][160] = 14'b11111111111111;
	assign font[9][160] = 14'b11111111111111;
	assign font[10][160] = 14'b11111111111111;
	assign font[11][160] = 14'b11111111111111;
	assign font[12][160] = 14'b11111111111111;
	assign font[13][160] = 14'b11111111111111;
	assign font[14][160] = 14'b11111111111111;
	assign font[15][160] = 14'b11111111111111;
	assign font[16][160] = 14'b11111111111111;
	assign font[17][160] = 14'b11111111111111;
	assign font[18][160] = 14'b11111111111111;
	assign font[19][160] = 14'b11111111111111;
	assign font[20][160] = 14'b11111111111111;
	assign font[21][160] = 14'b11111111111111;
	assign font[22][160] = 14'b11111111111111;
	assign font[23][160] = 14'b11111111111111;
	assign font[24][160] = 14'b11111111111111;
	assign font[25][160] = 14'b11111111111111;
	assign font[26][160] = 14'b11111111111111;
	assign font[27][160] = 14'b11111111111111;
	assign font[28][160] = 14'b11111111111111;
	assign font[29][160] = 14'b11111111111111;
	assign font[30][160] = 14'b11111111111111;
	assign font[31][160] = 14'b11111111111111;

	assign font[0][161] = 14'b11111111111111;
	assign font[1][161] = 14'b11111111111111;
	assign font[2][161] = 14'b11111111111111;
	assign font[3][161] = 14'b11111111111111;
	assign font[4][161] = 14'b11111111111111;
	assign font[5][161] = 14'b11111111111111;
	assign font[6][161] = 14'b11111111111111;
	assign font[7][161] = 14'b11111111111111;
	assign font[8][161] = 14'b11111111111111;
	assign font[9][161] = 14'b11111111111111;
	assign font[10][161] = 14'b11111111111111;
	assign font[11][161] = 14'b11111111111111;
	assign font[12][161] = 14'b11111111111111;
	assign font[13][161] = 14'b11111111111111;
	assign font[14][161] = 14'b11111111111111;
	assign font[15][161] = 14'b11111111111111;
	assign font[16][161] = 14'b11111111111111;
	assign font[17][161] = 14'b11111111111111;
	assign font[18][161] = 14'b11111111111111;
	assign font[19][161] = 14'b11111111111111;
	assign font[20][161] = 14'b11111111111111;
	assign font[21][161] = 14'b11111111111111;
	assign font[22][161] = 14'b11111111111111;
	assign font[23][161] = 14'b11111111111111;
	assign font[24][161] = 14'b11111111111111;
	assign font[25][161] = 14'b11111111111111;
	assign font[26][161] = 14'b11111111111111;
	assign font[27][161] = 14'b11111111111111;
	assign font[28][161] = 14'b11111111111111;
	assign font[29][161] = 14'b11111111111111;
	assign font[30][161] = 14'b11111111111111;
	assign font[31][161] = 14'b11111111111111;

	assign font[0][162] = 14'b11111111111111;
	assign font[1][162] = 14'b11111111111111;
	assign font[2][162] = 14'b11111111111111;
	assign font[3][162] = 14'b11111111111111;
	assign font[4][162] = 14'b11111111111111;
	assign font[5][162] = 14'b11111111111111;
	assign font[6][162] = 14'b11111111111111;
	assign font[7][162] = 14'b11111111111111;
	assign font[8][162] = 14'b11111111111111;
	assign font[9][162] = 14'b11111111111111;
	assign font[10][162] = 14'b11111111111111;
	assign font[11][162] = 14'b11111111111111;
	assign font[12][162] = 14'b11111111111111;
	assign font[13][162] = 14'b11111111111111;
	assign font[14][162] = 14'b11111111111111;
	assign font[15][162] = 14'b11111111111111;
	assign font[16][162] = 14'b11111111111111;
	assign font[17][162] = 14'b11111111111111;
	assign font[18][162] = 14'b11111111111111;
	assign font[19][162] = 14'b11111111111111;
	assign font[20][162] = 14'b11111111111111;
	assign font[21][162] = 14'b11111111111111;
	assign font[22][162] = 14'b11111111111111;
	assign font[23][162] = 14'b11111111111111;
	assign font[24][162] = 14'b11111111111111;
	assign font[25][162] = 14'b11111111111111;
	assign font[26][162] = 14'b11111111111111;
	assign font[27][162] = 14'b11111111111111;
	assign font[28][162] = 14'b11111111111111;
	assign font[29][162] = 14'b11111111111111;
	assign font[30][162] = 14'b11111111111111;
	assign font[31][162] = 14'b11111111111111;

	assign font[0][163] = 14'b11111111111111;
	assign font[1][163] = 14'b11111111111111;
	assign font[2][163] = 14'b11111111111111;
	assign font[3][163] = 14'b11111111111111;
	assign font[4][163] = 14'b11111111111111;
	assign font[5][163] = 14'b11111111111111;
	assign font[6][163] = 14'b11111111111111;
	assign font[7][163] = 14'b11111111111111;
	assign font[8][163] = 14'b11111111111111;
	assign font[9][163] = 14'b11111111111111;
	assign font[10][163] = 14'b11111111111111;
	assign font[11][163] = 14'b11111111111111;
	assign font[12][163] = 14'b11111111111111;
	assign font[13][163] = 14'b11111111111111;
	assign font[14][163] = 14'b11111111111111;
	assign font[15][163] = 14'b11111111111111;
	assign font[16][163] = 14'b11111111111111;
	assign font[17][163] = 14'b11111111111111;
	assign font[18][163] = 14'b11111111111111;
	assign font[19][163] = 14'b11111111111111;
	assign font[20][163] = 14'b11111111111111;
	assign font[21][163] = 14'b11111111111111;
	assign font[22][163] = 14'b11111111111111;
	assign font[23][163] = 14'b11111111111111;
	assign font[24][163] = 14'b11111111111111;
	assign font[25][163] = 14'b11111111111111;
	assign font[26][163] = 14'b11111111111111;
	assign font[27][163] = 14'b11111111111111;
	assign font[28][163] = 14'b11111111111111;
	assign font[29][163] = 14'b11111111111111;
	assign font[30][163] = 14'b11111111111111;
	assign font[31][163] = 14'b11111111111111;

	assign font[0][164] = 14'b11111111111111;
	assign font[1][164] = 14'b11111111111111;
	assign font[2][164] = 14'b11111111111111;
	assign font[3][164] = 14'b11111111111111;
	assign font[4][164] = 14'b11111111111111;
	assign font[5][164] = 14'b11111111111111;
	assign font[6][164] = 14'b11111111111111;
	assign font[7][164] = 14'b11111111111111;
	assign font[8][164] = 14'b11111111111111;
	assign font[9][164] = 14'b11111111111111;
	assign font[10][164] = 14'b11111111111111;
	assign font[11][164] = 14'b11111111111111;
	assign font[12][164] = 14'b11111111111111;
	assign font[13][164] = 14'b11111111111111;
	assign font[14][164] = 14'b11111111111111;
	assign font[15][164] = 14'b11111111111111;
	assign font[16][164] = 14'b11111111111111;
	assign font[17][164] = 14'b11111111111111;
	assign font[18][164] = 14'b11111111111111;
	assign font[19][164] = 14'b11111111111111;
	assign font[20][164] = 14'b11111111111111;
	assign font[21][164] = 14'b11111111111111;
	assign font[22][164] = 14'b11111111111111;
	assign font[23][164] = 14'b11111111111111;
	assign font[24][164] = 14'b11111111111111;
	assign font[25][164] = 14'b11111111111111;
	assign font[26][164] = 14'b11111111111111;
	assign font[27][164] = 14'b11111111111111;
	assign font[28][164] = 14'b11111111111111;
	assign font[29][164] = 14'b11111111111111;
	assign font[30][164] = 14'b11111111111111;
	assign font[31][164] = 14'b11111111111111;

	assign font[0][165] = 14'b11111111111111;
	assign font[1][165] = 14'b11111111111111;
	assign font[2][165] = 14'b11111111111111;
	assign font[3][165] = 14'b11111111111111;
	assign font[4][165] = 14'b11111111111111;
	assign font[5][165] = 14'b11111111111111;
	assign font[6][165] = 14'b11111111111111;
	assign font[7][165] = 14'b11111111111111;
	assign font[8][165] = 14'b11111111111111;
	assign font[9][165] = 14'b11111111111111;
	assign font[10][165] = 14'b11111111111111;
	assign font[11][165] = 14'b11111111111111;
	assign font[12][165] = 14'b11111111111111;
	assign font[13][165] = 14'b11111111111111;
	assign font[14][165] = 14'b11111111111111;
	assign font[15][165] = 14'b11111111111111;
	assign font[16][165] = 14'b11111111111111;
	assign font[17][165] = 14'b11111111111111;
	assign font[18][165] = 14'b11111111111111;
	assign font[19][165] = 14'b11111111111111;
	assign font[20][165] = 14'b11111111111111;
	assign font[21][165] = 14'b11111111111111;
	assign font[22][165] = 14'b11111111111111;
	assign font[23][165] = 14'b11111111111111;
	assign font[24][165] = 14'b11111111111111;
	assign font[25][165] = 14'b11111111111111;
	assign font[26][165] = 14'b11111111111111;
	assign font[27][165] = 14'b11111111111111;
	assign font[28][165] = 14'b11111111111111;
	assign font[29][165] = 14'b11111111111111;
	assign font[30][165] = 14'b11111111111111;
	assign font[31][165] = 14'b11111111111111;

	assign font[0][166] = 14'b11111111111111;
	assign font[1][166] = 14'b11111111111111;
	assign font[2][166] = 14'b11111111111111;
	assign font[3][166] = 14'b11111111111111;
	assign font[4][166] = 14'b11111111111111;
	assign font[5][166] = 14'b11111111111111;
	assign font[6][166] = 14'b11111111111111;
	assign font[7][166] = 14'b11111111111111;
	assign font[8][166] = 14'b11111111111111;
	assign font[9][166] = 14'b11111111111111;
	assign font[10][166] = 14'b11111111111111;
	assign font[11][166] = 14'b11111111111111;
	assign font[12][166] = 14'b11111111111111;
	assign font[13][166] = 14'b11111111111111;
	assign font[14][166] = 14'b11111111111111;
	assign font[15][166] = 14'b11111111111111;
	assign font[16][166] = 14'b11111111111111;
	assign font[17][166] = 14'b11111111111111;
	assign font[18][166] = 14'b11111111111111;
	assign font[19][166] = 14'b11111111111111;
	assign font[20][166] = 14'b11111111111111;
	assign font[21][166] = 14'b11111111111111;
	assign font[22][166] = 14'b11111111111111;
	assign font[23][166] = 14'b11111111111111;
	assign font[24][166] = 14'b11111111111111;
	assign font[25][166] = 14'b11111111111111;
	assign font[26][166] = 14'b11111111111111;
	assign font[27][166] = 14'b11111111111111;
	assign font[28][166] = 14'b11111111111111;
	assign font[29][166] = 14'b11111111111111;
	assign font[30][166] = 14'b11111111111111;
	assign font[31][166] = 14'b11111111111111;

	assign font[0][167] = 14'b11111111111111;
	assign font[1][167] = 14'b11111111111111;
	assign font[2][167] = 14'b11111111111111;
	assign font[3][167] = 14'b11111111111111;
	assign font[4][167] = 14'b11111111111111;
	assign font[5][167] = 14'b11111111111111;
	assign font[6][167] = 14'b11111111111111;
	assign font[7][167] = 14'b11111111111111;
	assign font[8][167] = 14'b11111111111111;
	assign font[9][167] = 14'b11111111111111;
	assign font[10][167] = 14'b11111111111111;
	assign font[11][167] = 14'b11111111111111;
	assign font[12][167] = 14'b11111111111111;
	assign font[13][167] = 14'b11111111111111;
	assign font[14][167] = 14'b11111111111111;
	assign font[15][167] = 14'b11111111111111;
	assign font[16][167] = 14'b11111111111111;
	assign font[17][167] = 14'b11111111111111;
	assign font[18][167] = 14'b11111111111111;
	assign font[19][167] = 14'b11111111111111;
	assign font[20][167] = 14'b11111111111111;
	assign font[21][167] = 14'b11111111111111;
	assign font[22][167] = 14'b11111111111111;
	assign font[23][167] = 14'b11111111111111;
	assign font[24][167] = 14'b11111111111111;
	assign font[25][167] = 14'b11111111111111;
	assign font[26][167] = 14'b11111111111111;
	assign font[27][167] = 14'b11111111111111;
	assign font[28][167] = 14'b11111111111111;
	assign font[29][167] = 14'b11111111111111;
	assign font[30][167] = 14'b11111111111111;
	assign font[31][167] = 14'b11111111111111;

	assign font[0][168] = 14'b11111111111111;
	assign font[1][168] = 14'b11111111111111;
	assign font[2][168] = 14'b11111111111111;
	assign font[3][168] = 14'b11111111111111;
	assign font[4][168] = 14'b11111111111111;
	assign font[5][168] = 14'b11111111111111;
	assign font[6][168] = 14'b11111111111111;
	assign font[7][168] = 14'b11111111111111;
	assign font[8][168] = 14'b11111111111111;
	assign font[9][168] = 14'b11111111111111;
	assign font[10][168] = 14'b11111111111111;
	assign font[11][168] = 14'b11111111111111;
	assign font[12][168] = 14'b11111111111111;
	assign font[13][168] = 14'b11111111111111;
	assign font[14][168] = 14'b11111111111111;
	assign font[15][168] = 14'b11111111111111;
	assign font[16][168] = 14'b11111111111111;
	assign font[17][168] = 14'b11111111111111;
	assign font[18][168] = 14'b11111111111111;
	assign font[19][168] = 14'b11111111111111;
	assign font[20][168] = 14'b11111111111111;
	assign font[21][168] = 14'b11111111111111;
	assign font[22][168] = 14'b11111111111111;
	assign font[23][168] = 14'b11111111111111;
	assign font[24][168] = 14'b11111111111111;
	assign font[25][168] = 14'b11111111111111;
	assign font[26][168] = 14'b11111111111111;
	assign font[27][168] = 14'b11111111111111;
	assign font[28][168] = 14'b11111111111111;
	assign font[29][168] = 14'b11111111111111;
	assign font[30][168] = 14'b11111111111111;
	assign font[31][168] = 14'b11111111111111;

	assign font[0][169] = 14'b11111111111111;
	assign font[1][169] = 14'b11111111111111;
	assign font[2][169] = 14'b11111111111111;
	assign font[3][169] = 14'b11111111111111;
	assign font[4][169] = 14'b11111111111111;
	assign font[5][169] = 14'b11111111111111;
	assign font[6][169] = 14'b11111111111111;
	assign font[7][169] = 14'b11111111111111;
	assign font[8][169] = 14'b11111111111111;
	assign font[9][169] = 14'b11111111111111;
	assign font[10][169] = 14'b11111111111111;
	assign font[11][169] = 14'b11111111111111;
	assign font[12][169] = 14'b11111111111111;
	assign font[13][169] = 14'b11111111111111;
	assign font[14][169] = 14'b11111111111111;
	assign font[15][169] = 14'b11111111111111;
	assign font[16][169] = 14'b11111111111111;
	assign font[17][169] = 14'b11111111111111;
	assign font[18][169] = 14'b11111111111111;
	assign font[19][169] = 14'b11111111111111;
	assign font[20][169] = 14'b11111111111111;
	assign font[21][169] = 14'b11111111111111;
	assign font[22][169] = 14'b11111111111111;
	assign font[23][169] = 14'b11111111111111;
	assign font[24][169] = 14'b11111111111111;
	assign font[25][169] = 14'b11111111111111;
	assign font[26][169] = 14'b11111111111111;
	assign font[27][169] = 14'b11111111111111;
	assign font[28][169] = 14'b11111111111111;
	assign font[29][169] = 14'b11111111111111;
	assign font[30][169] = 14'b11111111111111;
	assign font[31][169] = 14'b11111111111111;

	assign font[0][170] = 14'b11111111111111;
	assign font[1][170] = 14'b11111111111111;
	assign font[2][170] = 14'b11111111111111;
	assign font[3][170] = 14'b11111111111111;
	assign font[4][170] = 14'b11111111111111;
	assign font[5][170] = 14'b11111111111111;
	assign font[6][170] = 14'b11111111111111;
	assign font[7][170] = 14'b11111111111111;
	assign font[8][170] = 14'b11111111111111;
	assign font[9][170] = 14'b11111111111111;
	assign font[10][170] = 14'b11111111111111;
	assign font[11][170] = 14'b11111111111111;
	assign font[12][170] = 14'b11111111111111;
	assign font[13][170] = 14'b11111111111111;
	assign font[14][170] = 14'b11111111111111;
	assign font[15][170] = 14'b11111111111111;
	assign font[16][170] = 14'b11111111111111;
	assign font[17][170] = 14'b11111111111111;
	assign font[18][170] = 14'b11111111111111;
	assign font[19][170] = 14'b11111111111111;
	assign font[20][170] = 14'b11111111111111;
	assign font[21][170] = 14'b11111111111111;
	assign font[22][170] = 14'b11111111111111;
	assign font[23][170] = 14'b11111111111111;
	assign font[24][170] = 14'b11111111111111;
	assign font[25][170] = 14'b11111111111111;
	assign font[26][170] = 14'b11111111111111;
	assign font[27][170] = 14'b11111111111111;
	assign font[28][170] = 14'b11111111111111;
	assign font[29][170] = 14'b11111111111111;
	assign font[30][170] = 14'b11111111111111;
	assign font[31][170] = 14'b11111111111111;

	assign font[0][171] = 14'b11111111111111;
	assign font[1][171] = 14'b11111111111111;
	assign font[2][171] = 14'b11111111111111;
	assign font[3][171] = 14'b11111111111111;
	assign font[4][171] = 14'b11111111111111;
	assign font[5][171] = 14'b11111111111111;
	assign font[6][171] = 14'b11111111111111;
	assign font[7][171] = 14'b11111111111111;
	assign font[8][171] = 14'b11111111111111;
	assign font[9][171] = 14'b11111111111111;
	assign font[10][171] = 14'b11111111111111;
	assign font[11][171] = 14'b11111111111111;
	assign font[12][171] = 14'b11111111111111;
	assign font[13][171] = 14'b11111111111111;
	assign font[14][171] = 14'b11111111111111;
	assign font[15][171] = 14'b11111111111111;
	assign font[16][171] = 14'b11111111111111;
	assign font[17][171] = 14'b11111111111111;
	assign font[18][171] = 14'b11111111111111;
	assign font[19][171] = 14'b11111111111111;
	assign font[20][171] = 14'b11111111111111;
	assign font[21][171] = 14'b11111111111111;
	assign font[22][171] = 14'b11111111111111;
	assign font[23][171] = 14'b11111111111111;
	assign font[24][171] = 14'b11111111111111;
	assign font[25][171] = 14'b11111111111111;
	assign font[26][171] = 14'b11111111111111;
	assign font[27][171] = 14'b11111111111111;
	assign font[28][171] = 14'b11111111111111;
	assign font[29][171] = 14'b11111111111111;
	assign font[30][171] = 14'b11111111111111;
	assign font[31][171] = 14'b11111111111111;

	assign font[0][172] = 14'b11111111111111;
	assign font[1][172] = 14'b11111111111111;
	assign font[2][172] = 14'b11111111111111;
	assign font[3][172] = 14'b11111111111111;
	assign font[4][172] = 14'b11111111111111;
	assign font[5][172] = 14'b11111111111111;
	assign font[6][172] = 14'b11111111111111;
	assign font[7][172] = 14'b11111111111111;
	assign font[8][172] = 14'b11111111111111;
	assign font[9][172] = 14'b11111111111111;
	assign font[10][172] = 14'b11111111111111;
	assign font[11][172] = 14'b11111111111111;
	assign font[12][172] = 14'b11111111111111;
	assign font[13][172] = 14'b11111111111111;
	assign font[14][172] = 14'b11111111111111;
	assign font[15][172] = 14'b11111111111111;
	assign font[16][172] = 14'b11111111111111;
	assign font[17][172] = 14'b11111111111111;
	assign font[18][172] = 14'b11111111111111;
	assign font[19][172] = 14'b11111111111111;
	assign font[20][172] = 14'b11111111111111;
	assign font[21][172] = 14'b11111111111111;
	assign font[22][172] = 14'b11111111111111;
	assign font[23][172] = 14'b11111111111111;
	assign font[24][172] = 14'b11111111111111;
	assign font[25][172] = 14'b11111111111111;
	assign font[26][172] = 14'b11111111111111;
	assign font[27][172] = 14'b11111111111111;
	assign font[28][172] = 14'b11111111111111;
	assign font[29][172] = 14'b11111111111111;
	assign font[30][172] = 14'b11111111111111;
	assign font[31][172] = 14'b11111111111111;

	assign font[0][173] = 14'b11111111111111;
	assign font[1][173] = 14'b11111111111111;
	assign font[2][173] = 14'b11111111111111;
	assign font[3][173] = 14'b11111111111111;
	assign font[4][173] = 14'b11111111111111;
	assign font[5][173] = 14'b11111111111111;
	assign font[6][173] = 14'b11111111111111;
	assign font[7][173] = 14'b11111111111111;
	assign font[8][173] = 14'b11111111111111;
	assign font[9][173] = 14'b11111111111111;
	assign font[10][173] = 14'b11111111111111;
	assign font[11][173] = 14'b11111111111111;
	assign font[12][173] = 14'b11111111111111;
	assign font[13][173] = 14'b11111111111111;
	assign font[14][173] = 14'b11111111111111;
	assign font[15][173] = 14'b11111111111111;
	assign font[16][173] = 14'b11111111111111;
	assign font[17][173] = 14'b11111111111111;
	assign font[18][173] = 14'b11111111111111;
	assign font[19][173] = 14'b11111111111111;
	assign font[20][173] = 14'b11111111111111;
	assign font[21][173] = 14'b11111111111111;
	assign font[22][173] = 14'b11111111111111;
	assign font[23][173] = 14'b11111111111111;
	assign font[24][173] = 14'b11111111111111;
	assign font[25][173] = 14'b11111111111111;
	assign font[26][173] = 14'b11111111111111;
	assign font[27][173] = 14'b11111111111111;
	assign font[28][173] = 14'b11111111111111;
	assign font[29][173] = 14'b11111111111111;
	assign font[30][173] = 14'b11111111111111;
	assign font[31][173] = 14'b11111111111111;

	assign font[0][174] = 14'b11111111111111;
	assign font[1][174] = 14'b11111111111111;
	assign font[2][174] = 14'b11111111111111;
	assign font[3][174] = 14'b11111111111111;
	assign font[4][174] = 14'b11111111111111;
	assign font[5][174] = 14'b11111111111111;
	assign font[6][174] = 14'b11111111111111;
	assign font[7][174] = 14'b11111111111111;
	assign font[8][174] = 14'b11111111111111;
	assign font[9][174] = 14'b11111111111111;
	assign font[10][174] = 14'b11111111111111;
	assign font[11][174] = 14'b11111111111111;
	assign font[12][174] = 14'b11111111111111;
	assign font[13][174] = 14'b11111111111111;
	assign font[14][174] = 14'b11111111111111;
	assign font[15][174] = 14'b11111111111111;
	assign font[16][174] = 14'b11111111111111;
	assign font[17][174] = 14'b11111111111111;
	assign font[18][174] = 14'b11111111111111;
	assign font[19][174] = 14'b11111111111111;
	assign font[20][174] = 14'b11111111111111;
	assign font[21][174] = 14'b11111111111111;
	assign font[22][174] = 14'b11111111111111;
	assign font[23][174] = 14'b11111111111111;
	assign font[24][174] = 14'b11111111111111;
	assign font[25][174] = 14'b11111111111111;
	assign font[26][174] = 14'b11111111111111;
	assign font[27][174] = 14'b11111111111111;
	assign font[28][174] = 14'b11111111111111;
	assign font[29][174] = 14'b11111111111111;
	assign font[30][174] = 14'b11111111111111;
	assign font[31][174] = 14'b11111111111111;

	assign font[0][175] = 14'b11111111111111;
	assign font[1][175] = 14'b11111111111111;
	assign font[2][175] = 14'b11111111111111;
	assign font[3][175] = 14'b11111111111111;
	assign font[4][175] = 14'b11111111111111;
	assign font[5][175] = 14'b11111111111111;
	assign font[6][175] = 14'b11111111111111;
	assign font[7][175] = 14'b11111111111111;
	assign font[8][175] = 14'b11111111111111;
	assign font[9][175] = 14'b11111111111111;
	assign font[10][175] = 14'b11111111111111;
	assign font[11][175] = 14'b11111111111111;
	assign font[12][175] = 14'b11111111111111;
	assign font[13][175] = 14'b11111111111111;
	assign font[14][175] = 14'b11111111111111;
	assign font[15][175] = 14'b11111111111111;
	assign font[16][175] = 14'b11111111111111;
	assign font[17][175] = 14'b11111111111111;
	assign font[18][175] = 14'b11111111111111;
	assign font[19][175] = 14'b11111111111111;
	assign font[20][175] = 14'b11111111111111;
	assign font[21][175] = 14'b11111111111111;
	assign font[22][175] = 14'b11111111111111;
	assign font[23][175] = 14'b11111111111111;
	assign font[24][175] = 14'b11111111111111;
	assign font[25][175] = 14'b11111111111111;
	assign font[26][175] = 14'b11111111111111;
	assign font[27][175] = 14'b11111111111111;
	assign font[28][175] = 14'b11111111111111;
	assign font[29][175] = 14'b11111111111111;
	assign font[30][175] = 14'b11111111111111;
	assign font[31][175] = 14'b11111111111111;

	assign font[0][176] = 14'b11111111111111;
	assign font[1][176] = 14'b11111111111111;
	assign font[2][176] = 14'b11111111111111;
	assign font[3][176] = 14'b11111111111111;
	assign font[4][176] = 14'b11111111111111;
	assign font[5][176] = 14'b11111111111111;
	assign font[6][176] = 14'b11111111111111;
	assign font[7][176] = 14'b11111111111111;
	assign font[8][176] = 14'b11111111111111;
	assign font[9][176] = 14'b11111111111111;
	assign font[10][176] = 14'b11111111111111;
	assign font[11][176] = 14'b11111111111111;
	assign font[12][176] = 14'b11111111111111;
	assign font[13][176] = 14'b11111111111111;
	assign font[14][176] = 14'b11111111111111;
	assign font[15][176] = 14'b11111111111111;
	assign font[16][176] = 14'b11111111111111;
	assign font[17][176] = 14'b11111111111111;
	assign font[18][176] = 14'b11111111111111;
	assign font[19][176] = 14'b11111111111111;
	assign font[20][176] = 14'b11111111111111;
	assign font[21][176] = 14'b11111111111111;
	assign font[22][176] = 14'b11111111111111;
	assign font[23][176] = 14'b11111111111111;
	assign font[24][176] = 14'b11111111111111;
	assign font[25][176] = 14'b11111111111111;
	assign font[26][176] = 14'b11111111111111;
	assign font[27][176] = 14'b11111111111111;
	assign font[28][176] = 14'b11111111111111;
	assign font[29][176] = 14'b11111111111111;
	assign font[30][176] = 14'b11111111111111;
	assign font[31][176] = 14'b11111111111111;

	assign font[0][177] = 14'b11111111111111;
	assign font[1][177] = 14'b11111111111111;
	assign font[2][177] = 14'b11111111111111;
	assign font[3][177] = 14'b11111111111111;
	assign font[4][177] = 14'b11111111111111;
	assign font[5][177] = 14'b11111111111111;
	assign font[6][177] = 14'b11111111111111;
	assign font[7][177] = 14'b11111111111111;
	assign font[8][177] = 14'b11111111111111;
	assign font[9][177] = 14'b11111111111111;
	assign font[10][177] = 14'b11111111111111;
	assign font[11][177] = 14'b11111111111111;
	assign font[12][177] = 14'b11111111111111;
	assign font[13][177] = 14'b11111111111111;
	assign font[14][177] = 14'b11111111111111;
	assign font[15][177] = 14'b11111111111111;
	assign font[16][177] = 14'b11111111111111;
	assign font[17][177] = 14'b11111111111111;
	assign font[18][177] = 14'b11111111111111;
	assign font[19][177] = 14'b11111111111111;
	assign font[20][177] = 14'b11111111111111;
	assign font[21][177] = 14'b11111111111111;
	assign font[22][177] = 14'b11111111111111;
	assign font[23][177] = 14'b11111111111111;
	assign font[24][177] = 14'b11111111111111;
	assign font[25][177] = 14'b11111111111111;
	assign font[26][177] = 14'b11111111111111;
	assign font[27][177] = 14'b11111111111111;
	assign font[28][177] = 14'b11111111111111;
	assign font[29][177] = 14'b11111111111111;
	assign font[30][177] = 14'b11111111111111;
	assign font[31][177] = 14'b11111111111111;

	assign font[0][178] = 14'b11111111111111;
	assign font[1][178] = 14'b11111111111111;
	assign font[2][178] = 14'b11111111111111;
	assign font[3][178] = 14'b11111111111111;
	assign font[4][178] = 14'b11111111111111;
	assign font[5][178] = 14'b11111111111111;
	assign font[6][178] = 14'b11111111111111;
	assign font[7][178] = 14'b11111111111111;
	assign font[8][178] = 14'b11111111111111;
	assign font[9][178] = 14'b11111111111111;
	assign font[10][178] = 14'b11111111111111;
	assign font[11][178] = 14'b11111111111111;
	assign font[12][178] = 14'b11111111111111;
	assign font[13][178] = 14'b11111111111111;
	assign font[14][178] = 14'b11111111111111;
	assign font[15][178] = 14'b11111111111111;
	assign font[16][178] = 14'b11111111111111;
	assign font[17][178] = 14'b11111111111111;
	assign font[18][178] = 14'b11111111111111;
	assign font[19][178] = 14'b11111111111111;
	assign font[20][178] = 14'b11111111111111;
	assign font[21][178] = 14'b11111111111111;
	assign font[22][178] = 14'b11111111111111;
	assign font[23][178] = 14'b11111111111111;
	assign font[24][178] = 14'b11111111111111;
	assign font[25][178] = 14'b11111111111111;
	assign font[26][178] = 14'b11111111111111;
	assign font[27][178] = 14'b11111111111111;
	assign font[28][178] = 14'b11111111111111;
	assign font[29][178] = 14'b11111111111111;
	assign font[30][178] = 14'b11111111111111;
	assign font[31][178] = 14'b11111111111111;

	assign font[0][179] = 14'b11111111111111;
	assign font[1][179] = 14'b11111111111111;
	assign font[2][179] = 14'b11111111111111;
	assign font[3][179] = 14'b11111111111111;
	assign font[4][179] = 14'b11111111111111;
	assign font[5][179] = 14'b11111111111111;
	assign font[6][179] = 14'b11111111111111;
	assign font[7][179] = 14'b11111111111111;
	assign font[8][179] = 14'b11111111111111;
	assign font[9][179] = 14'b11111111111111;
	assign font[10][179] = 14'b11111111111111;
	assign font[11][179] = 14'b11111111111111;
	assign font[12][179] = 14'b11111111111111;
	assign font[13][179] = 14'b11111111111111;
	assign font[14][179] = 14'b11111111111111;
	assign font[15][179] = 14'b11111111111111;
	assign font[16][179] = 14'b11111111111111;
	assign font[17][179] = 14'b11111111111111;
	assign font[18][179] = 14'b11111111111111;
	assign font[19][179] = 14'b11111111111111;
	assign font[20][179] = 14'b11111111111111;
	assign font[21][179] = 14'b11111111111111;
	assign font[22][179] = 14'b11111111111111;
	assign font[23][179] = 14'b11111111111111;
	assign font[24][179] = 14'b11111111111111;
	assign font[25][179] = 14'b11111111111111;
	assign font[26][179] = 14'b11111111111111;
	assign font[27][179] = 14'b11111111111111;
	assign font[28][179] = 14'b11111111111111;
	assign font[29][179] = 14'b11111111111111;
	assign font[30][179] = 14'b11111111111111;
	assign font[31][179] = 14'b11111111111111;

	assign font[0][180] = 14'b11111111111111;
	assign font[1][180] = 14'b11111111111111;
	assign font[2][180] = 14'b11111111111111;
	assign font[3][180] = 14'b11111111111111;
	assign font[4][180] = 14'b11111111111111;
	assign font[5][180] = 14'b11111111111111;
	assign font[6][180] = 14'b11111111111111;
	assign font[7][180] = 14'b11111111111111;
	assign font[8][180] = 14'b11111111111111;
	assign font[9][180] = 14'b11111111111111;
	assign font[10][180] = 14'b11111111111111;
	assign font[11][180] = 14'b11111111111111;
	assign font[12][180] = 14'b11111111111111;
	assign font[13][180] = 14'b11111111111111;
	assign font[14][180] = 14'b11111111111111;
	assign font[15][180] = 14'b11111111111111;
	assign font[16][180] = 14'b11111111111111;
	assign font[17][180] = 14'b11111111111111;
	assign font[18][180] = 14'b11111111111111;
	assign font[19][180] = 14'b11111111111111;
	assign font[20][180] = 14'b11111111111111;
	assign font[21][180] = 14'b11111111111111;
	assign font[22][180] = 14'b11111111111111;
	assign font[23][180] = 14'b11111111111111;
	assign font[24][180] = 14'b11111111111111;
	assign font[25][180] = 14'b11111111111111;
	assign font[26][180] = 14'b11111111111111;
	assign font[27][180] = 14'b11111111111111;
	assign font[28][180] = 14'b11111111111111;
	assign font[29][180] = 14'b11111111111111;
	assign font[30][180] = 14'b11111111111111;
	assign font[31][180] = 14'b11111111111111;

	assign font[0][181] = 14'b11111111111111;
	assign font[1][181] = 14'b11111111111111;
	assign font[2][181] = 14'b11111111111111;
	assign font[3][181] = 14'b11111111111111;
	assign font[4][181] = 14'b11111111111111;
	assign font[5][181] = 14'b11111111111111;
	assign font[6][181] = 14'b11111111111111;
	assign font[7][181] = 14'b11111111111111;
	assign font[8][181] = 14'b11111111111111;
	assign font[9][181] = 14'b11111111111111;
	assign font[10][181] = 14'b11111111111111;
	assign font[11][181] = 14'b11111111111111;
	assign font[12][181] = 14'b11111111111111;
	assign font[13][181] = 14'b11111111111111;
	assign font[14][181] = 14'b11111111111111;
	assign font[15][181] = 14'b11111111111111;
	assign font[16][181] = 14'b11111111111111;
	assign font[17][181] = 14'b11111111111111;
	assign font[18][181] = 14'b11111111111111;
	assign font[19][181] = 14'b11111111111111;
	assign font[20][181] = 14'b11111111111111;
	assign font[21][181] = 14'b11111111111111;
	assign font[22][181] = 14'b11111111111111;
	assign font[23][181] = 14'b11111111111111;
	assign font[24][181] = 14'b11111111111111;
	assign font[25][181] = 14'b11111111111111;
	assign font[26][181] = 14'b11111111111111;
	assign font[27][181] = 14'b11111111111111;
	assign font[28][181] = 14'b11111111111111;
	assign font[29][181] = 14'b11111111111111;
	assign font[30][181] = 14'b11111111111111;
	assign font[31][181] = 14'b11111111111111;

	assign font[0][182] = 14'b11111111111111;
	assign font[1][182] = 14'b11111111111111;
	assign font[2][182] = 14'b11111111111111;
	assign font[3][182] = 14'b11111111111111;
	assign font[4][182] = 14'b11111111111111;
	assign font[5][182] = 14'b11111111111111;
	assign font[6][182] = 14'b11111111111111;
	assign font[7][182] = 14'b11111111111111;
	assign font[8][182] = 14'b11111111111111;
	assign font[9][182] = 14'b11111111111111;
	assign font[10][182] = 14'b11111111111111;
	assign font[11][182] = 14'b11111111111111;
	assign font[12][182] = 14'b11111111111111;
	assign font[13][182] = 14'b11111111111111;
	assign font[14][182] = 14'b11111111111111;
	assign font[15][182] = 14'b11111111111111;
	assign font[16][182] = 14'b11111111111111;
	assign font[17][182] = 14'b11111111111111;
	assign font[18][182] = 14'b11111111111111;
	assign font[19][182] = 14'b11111111111111;
	assign font[20][182] = 14'b11111111111111;
	assign font[21][182] = 14'b11111111111111;
	assign font[22][182] = 14'b11111111111111;
	assign font[23][182] = 14'b11111111111111;
	assign font[24][182] = 14'b11111111111111;
	assign font[25][182] = 14'b11111111111111;
	assign font[26][182] = 14'b11111111111111;
	assign font[27][182] = 14'b11111111111111;
	assign font[28][182] = 14'b11111111111111;
	assign font[29][182] = 14'b11111111111111;
	assign font[30][182] = 14'b11111111111111;
	assign font[31][182] = 14'b11111111111111;

	assign font[0][183] = 14'b11111111111111;
	assign font[1][183] = 14'b11111111111111;
	assign font[2][183] = 14'b11111111111111;
	assign font[3][183] = 14'b11111111111111;
	assign font[4][183] = 14'b11111111111111;
	assign font[5][183] = 14'b11111111111111;
	assign font[6][183] = 14'b11111111111111;
	assign font[7][183] = 14'b11111111111111;
	assign font[8][183] = 14'b11111111111111;
	assign font[9][183] = 14'b11111111111111;
	assign font[10][183] = 14'b11111111111111;
	assign font[11][183] = 14'b11111111111111;
	assign font[12][183] = 14'b11111111111111;
	assign font[13][183] = 14'b11111111111111;
	assign font[14][183] = 14'b11111111111111;
	assign font[15][183] = 14'b11111111111111;
	assign font[16][183] = 14'b11111111111111;
	assign font[17][183] = 14'b11111111111111;
	assign font[18][183] = 14'b11111111111111;
	assign font[19][183] = 14'b11111111111111;
	assign font[20][183] = 14'b11111111111111;
	assign font[21][183] = 14'b11111111111111;
	assign font[22][183] = 14'b11111111111111;
	assign font[23][183] = 14'b11111111111111;
	assign font[24][183] = 14'b11111111111111;
	assign font[25][183] = 14'b11111111111111;
	assign font[26][183] = 14'b11111111111111;
	assign font[27][183] = 14'b11111111111111;
	assign font[28][183] = 14'b11111111111111;
	assign font[29][183] = 14'b11111111111111;
	assign font[30][183] = 14'b11111111111111;
	assign font[31][183] = 14'b11111111111111;

	assign font[0][184] = 14'b11111111111111;
	assign font[1][184] = 14'b11111111111111;
	assign font[2][184] = 14'b11111111111111;
	assign font[3][184] = 14'b11111111111111;
	assign font[4][184] = 14'b11111111111111;
	assign font[5][184] = 14'b11111111111111;
	assign font[6][184] = 14'b11111111111111;
	assign font[7][184] = 14'b11111111111111;
	assign font[8][184] = 14'b11111111111111;
	assign font[9][184] = 14'b11111111111111;
	assign font[10][184] = 14'b11111111111111;
	assign font[11][184] = 14'b11111111111111;
	assign font[12][184] = 14'b11111111111111;
	assign font[13][184] = 14'b11111111111111;
	assign font[14][184] = 14'b11111111111111;
	assign font[15][184] = 14'b11111111111111;
	assign font[16][184] = 14'b11111111111111;
	assign font[17][184] = 14'b11111111111111;
	assign font[18][184] = 14'b11111111111111;
	assign font[19][184] = 14'b11111111111111;
	assign font[20][184] = 14'b11111111111111;
	assign font[21][184] = 14'b11111111111111;
	assign font[22][184] = 14'b11111111111111;
	assign font[23][184] = 14'b11111111111111;
	assign font[24][184] = 14'b11111111111111;
	assign font[25][184] = 14'b11111111111111;
	assign font[26][184] = 14'b11111111111111;
	assign font[27][184] = 14'b11111111111111;
	assign font[28][184] = 14'b11111111111111;
	assign font[29][184] = 14'b11111111111111;
	assign font[30][184] = 14'b11111111111111;
	assign font[31][184] = 14'b11111111111111;

	assign font[0][185] = 14'b11111111111111;
	assign font[1][185] = 14'b11111111111111;
	assign font[2][185] = 14'b11111111111111;
	assign font[3][185] = 14'b11111111111111;
	assign font[4][185] = 14'b11111111111111;
	assign font[5][185] = 14'b11111111111111;
	assign font[6][185] = 14'b11111111111111;
	assign font[7][185] = 14'b11111111111111;
	assign font[8][185] = 14'b11111111111111;
	assign font[9][185] = 14'b11111111111111;
	assign font[10][185] = 14'b11111111111111;
	assign font[11][185] = 14'b11111111111111;
	assign font[12][185] = 14'b11111111111111;
	assign font[13][185] = 14'b11111111111111;
	assign font[14][185] = 14'b11111111111111;
	assign font[15][185] = 14'b11111111111111;
	assign font[16][185] = 14'b11111111111111;
	assign font[17][185] = 14'b11111111111111;
	assign font[18][185] = 14'b11111111111111;
	assign font[19][185] = 14'b11111111111111;
	assign font[20][185] = 14'b11111111111111;
	assign font[21][185] = 14'b11111111111111;
	assign font[22][185] = 14'b11111111111111;
	assign font[23][185] = 14'b11111111111111;
	assign font[24][185] = 14'b11111111111111;
	assign font[25][185] = 14'b11111111111111;
	assign font[26][185] = 14'b11111111111111;
	assign font[27][185] = 14'b11111111111111;
	assign font[28][185] = 14'b11111111111111;
	assign font[29][185] = 14'b11111111111111;
	assign font[30][185] = 14'b11111111111111;
	assign font[31][185] = 14'b11111111111111;

	assign font[0][186] = 14'b11111111111111;
	assign font[1][186] = 14'b11111111111111;
	assign font[2][186] = 14'b11111111111111;
	assign font[3][186] = 14'b11111111111111;
	assign font[4][186] = 14'b11111111111111;
	assign font[5][186] = 14'b11111111111111;
	assign font[6][186] = 14'b11111111111111;
	assign font[7][186] = 14'b11111111111111;
	assign font[8][186] = 14'b11111111111111;
	assign font[9][186] = 14'b11111111111111;
	assign font[10][186] = 14'b11111111111111;
	assign font[11][186] = 14'b11111111111111;
	assign font[12][186] = 14'b11111111111111;
	assign font[13][186] = 14'b11111111111111;
	assign font[14][186] = 14'b11111111111111;
	assign font[15][186] = 14'b11111111111111;
	assign font[16][186] = 14'b11111111111111;
	assign font[17][186] = 14'b11111111111111;
	assign font[18][186] = 14'b11111111111111;
	assign font[19][186] = 14'b11111111111111;
	assign font[20][186] = 14'b11111111111111;
	assign font[21][186] = 14'b11111111111111;
	assign font[22][186] = 14'b11111111111111;
	assign font[23][186] = 14'b11111111111111;
	assign font[24][186] = 14'b11111111111111;
	assign font[25][186] = 14'b11111111111111;
	assign font[26][186] = 14'b11111111111111;
	assign font[27][186] = 14'b11111111111111;
	assign font[28][186] = 14'b11111111111111;
	assign font[29][186] = 14'b11111111111111;
	assign font[30][186] = 14'b11111111111111;
	assign font[31][186] = 14'b11111111111111;

	assign font[0][187] = 14'b11111111111111;
	assign font[1][187] = 14'b11111111111111;
	assign font[2][187] = 14'b11111111111111;
	assign font[3][187] = 14'b11111111111111;
	assign font[4][187] = 14'b11111111111111;
	assign font[5][187] = 14'b11111111111111;
	assign font[6][187] = 14'b11111111111111;
	assign font[7][187] = 14'b11111111111111;
	assign font[8][187] = 14'b11111111111111;
	assign font[9][187] = 14'b11111111111111;
	assign font[10][187] = 14'b11111111111111;
	assign font[11][187] = 14'b11111111111111;
	assign font[12][187] = 14'b11111111111111;
	assign font[13][187] = 14'b11111111111111;
	assign font[14][187] = 14'b11111111111111;
	assign font[15][187] = 14'b11111111111111;
	assign font[16][187] = 14'b11111111111111;
	assign font[17][187] = 14'b11111111111111;
	assign font[18][187] = 14'b11111111111111;
	assign font[19][187] = 14'b11111111111111;
	assign font[20][187] = 14'b11111111111111;
	assign font[21][187] = 14'b11111111111111;
	assign font[22][187] = 14'b11111111111111;
	assign font[23][187] = 14'b11111111111111;
	assign font[24][187] = 14'b11111111111111;
	assign font[25][187] = 14'b11111111111111;
	assign font[26][187] = 14'b11111111111111;
	assign font[27][187] = 14'b11111111111111;
	assign font[28][187] = 14'b11111111111111;
	assign font[29][187] = 14'b11111111111111;
	assign font[30][187] = 14'b11111111111111;
	assign font[31][187] = 14'b11111111111111;

	assign font[0][188] = 14'b11111111111111;
	assign font[1][188] = 14'b11111111111111;
	assign font[2][188] = 14'b11111111111111;
	assign font[3][188] = 14'b11111111111111;
	assign font[4][188] = 14'b11111111111111;
	assign font[5][188] = 14'b11111111111111;
	assign font[6][188] = 14'b11111111111111;
	assign font[7][188] = 14'b11111111111111;
	assign font[8][188] = 14'b11111111111111;
	assign font[9][188] = 14'b11111111111111;
	assign font[10][188] = 14'b11111111111111;
	assign font[11][188] = 14'b11111111111111;
	assign font[12][188] = 14'b11111111111111;
	assign font[13][188] = 14'b11111111111111;
	assign font[14][188] = 14'b11111111111111;
	assign font[15][188] = 14'b11111111111111;
	assign font[16][188] = 14'b11111111111111;
	assign font[17][188] = 14'b11111111111111;
	assign font[18][188] = 14'b11111111111111;
	assign font[19][188] = 14'b11111111111111;
	assign font[20][188] = 14'b11111111111111;
	assign font[21][188] = 14'b11111111111111;
	assign font[22][188] = 14'b11111111111111;
	assign font[23][188] = 14'b11111111111111;
	assign font[24][188] = 14'b11111111111111;
	assign font[25][188] = 14'b11111111111111;
	assign font[26][188] = 14'b11111111111111;
	assign font[27][188] = 14'b11111111111111;
	assign font[28][188] = 14'b11111111111111;
	assign font[29][188] = 14'b11111111111111;
	assign font[30][188] = 14'b11111111111111;
	assign font[31][188] = 14'b11111111111111;

	assign font[0][189] = 14'b11111111111111;
	assign font[1][189] = 14'b11111111111111;
	assign font[2][189] = 14'b11111111111111;
	assign font[3][189] = 14'b11111111111111;
	assign font[4][189] = 14'b11111111111111;
	assign font[5][189] = 14'b11111111111111;
	assign font[6][189] = 14'b11111111111111;
	assign font[7][189] = 14'b11111111111111;
	assign font[8][189] = 14'b11111111111111;
	assign font[9][189] = 14'b11111111111111;
	assign font[10][189] = 14'b11111111111111;
	assign font[11][189] = 14'b11111111111111;
	assign font[12][189] = 14'b11111111111111;
	assign font[13][189] = 14'b11111111111111;
	assign font[14][189] = 14'b11111111111111;
	assign font[15][189] = 14'b11111111111111;
	assign font[16][189] = 14'b11111111111111;
	assign font[17][189] = 14'b11111111111111;
	assign font[18][189] = 14'b11111111111111;
	assign font[19][189] = 14'b11111111111111;
	assign font[20][189] = 14'b11111111111111;
	assign font[21][189] = 14'b11111111111111;
	assign font[22][189] = 14'b11111111111111;
	assign font[23][189] = 14'b11111111111111;
	assign font[24][189] = 14'b11111111111111;
	assign font[25][189] = 14'b11111111111111;
	assign font[26][189] = 14'b11111111111111;
	assign font[27][189] = 14'b11111111111111;
	assign font[28][189] = 14'b11111111111111;
	assign font[29][189] = 14'b11111111111111;
	assign font[30][189] = 14'b11111111111111;
	assign font[31][189] = 14'b11111111111111;

	assign font[0][190] = 14'b11111111111111;
	assign font[1][190] = 14'b11111111111111;
	assign font[2][190] = 14'b11111111111111;
	assign font[3][190] = 14'b11111111111111;
	assign font[4][190] = 14'b11111111111111;
	assign font[5][190] = 14'b11111111111111;
	assign font[6][190] = 14'b11111111111111;
	assign font[7][190] = 14'b11111111111111;
	assign font[8][190] = 14'b11111111111111;
	assign font[9][190] = 14'b11111111111111;
	assign font[10][190] = 14'b11111111111111;
	assign font[11][190] = 14'b11111111111111;
	assign font[12][190] = 14'b11111111111111;
	assign font[13][190] = 14'b11111111111111;
	assign font[14][190] = 14'b11111111111111;
	assign font[15][190] = 14'b11111111111111;
	assign font[16][190] = 14'b11111111111111;
	assign font[17][190] = 14'b11111111111111;
	assign font[18][190] = 14'b11111111111111;
	assign font[19][190] = 14'b11111111111111;
	assign font[20][190] = 14'b11111111111111;
	assign font[21][190] = 14'b11111111111111;
	assign font[22][190] = 14'b11111111111111;
	assign font[23][190] = 14'b11111111111111;
	assign font[24][190] = 14'b11111111111111;
	assign font[25][190] = 14'b11111111111111;
	assign font[26][190] = 14'b11111111111111;
	assign font[27][190] = 14'b11111111111111;
	assign font[28][190] = 14'b11111111111111;
	assign font[29][190] = 14'b11111111111111;
	assign font[30][190] = 14'b11111111111111;
	assign font[31][190] = 14'b11111111111111;

	assign font[0][191] = 14'b11111111111111;
	assign font[1][191] = 14'b11111111111111;
	assign font[2][191] = 14'b11111111111111;
	assign font[3][191] = 14'b11111111111111;
	assign font[4][191] = 14'b11111111111111;
	assign font[5][191] = 14'b11111111111111;
	assign font[6][191] = 14'b11111111111111;
	assign font[7][191] = 14'b11111111111111;
	assign font[8][191] = 14'b11111111111111;
	assign font[9][191] = 14'b11111111111111;
	assign font[10][191] = 14'b11111111111111;
	assign font[11][191] = 14'b11111111111111;
	assign font[12][191] = 14'b11111111111111;
	assign font[13][191] = 14'b11111111111111;
	assign font[14][191] = 14'b11111111111111;
	assign font[15][191] = 14'b11111111111111;
	assign font[16][191] = 14'b11111111111111;
	assign font[17][191] = 14'b11111111111111;
	assign font[18][191] = 14'b11111111111111;
	assign font[19][191] = 14'b11111111111111;
	assign font[20][191] = 14'b11111111111111;
	assign font[21][191] = 14'b11111111111111;
	assign font[22][191] = 14'b11111111111111;
	assign font[23][191] = 14'b11111111111111;
	assign font[24][191] = 14'b11111111111111;
	assign font[25][191] = 14'b11111111111111;
	assign font[26][191] = 14'b11111111111111;
	assign font[27][191] = 14'b11111111111111;
	assign font[28][191] = 14'b11111111111111;
	assign font[29][191] = 14'b11111111111111;
	assign font[30][191] = 14'b11111111111111;
	assign font[31][191] = 14'b11111111111111;

	assign font[0][192] = 14'b11111111111111;
	assign font[1][192] = 14'b11111111111111;
	assign font[2][192] = 14'b11111111111111;
	assign font[3][192] = 14'b11111111111111;
	assign font[4][192] = 14'b11111111111111;
	assign font[5][192] = 14'b11111111111111;
	assign font[6][192] = 14'b11111111111111;
	assign font[7][192] = 14'b11111111111111;
	assign font[8][192] = 14'b11111111111111;
	assign font[9][192] = 14'b11111111111111;
	assign font[10][192] = 14'b11111111111111;
	assign font[11][192] = 14'b11111111111111;
	assign font[12][192] = 14'b11111111111111;
	assign font[13][192] = 14'b11111111111111;
	assign font[14][192] = 14'b11111111111111;
	assign font[15][192] = 14'b11111111111111;
	assign font[16][192] = 14'b11111111111111;
	assign font[17][192] = 14'b11111111111111;
	assign font[18][192] = 14'b11111111111111;
	assign font[19][192] = 14'b11111111111111;
	assign font[20][192] = 14'b11111111111111;
	assign font[21][192] = 14'b11111111111111;
	assign font[22][192] = 14'b11111111111111;
	assign font[23][192] = 14'b11111111111111;
	assign font[24][192] = 14'b11111111111111;
	assign font[25][192] = 14'b11111111111111;
	assign font[26][192] = 14'b11111111111111;
	assign font[27][192] = 14'b11111111111111;
	assign font[28][192] = 14'b11111111111111;
	assign font[29][192] = 14'b11111111111111;
	assign font[30][192] = 14'b11111111111111;
	assign font[31][192] = 14'b11111111111111;

	assign font[0][193] = 14'b11111111111111;
	assign font[1][193] = 14'b11111111111111;
	assign font[2][193] = 14'b11111111111111;
	assign font[3][193] = 14'b11111111111111;
	assign font[4][193] = 14'b11111111111111;
	assign font[5][193] = 14'b11111111111111;
	assign font[6][193] = 14'b11111111111111;
	assign font[7][193] = 14'b11111111111111;
	assign font[8][193] = 14'b11111111111111;
	assign font[9][193] = 14'b11111111111111;
	assign font[10][193] = 14'b11111111111111;
	assign font[11][193] = 14'b11111111111111;
	assign font[12][193] = 14'b11111111111111;
	assign font[13][193] = 14'b11111111111111;
	assign font[14][193] = 14'b11111111111111;
	assign font[15][193] = 14'b11111111111111;
	assign font[16][193] = 14'b11111111111111;
	assign font[17][193] = 14'b11111111111111;
	assign font[18][193] = 14'b11111111111111;
	assign font[19][193] = 14'b11111111111111;
	assign font[20][193] = 14'b11111111111111;
	assign font[21][193] = 14'b11111111111111;
	assign font[22][193] = 14'b11111111111111;
	assign font[23][193] = 14'b11111111111111;
	assign font[24][193] = 14'b11111111111111;
	assign font[25][193] = 14'b11111111111111;
	assign font[26][193] = 14'b11111111111111;
	assign font[27][193] = 14'b11111111111111;
	assign font[28][193] = 14'b11111111111111;
	assign font[29][193] = 14'b11111111111111;
	assign font[30][193] = 14'b11111111111111;
	assign font[31][193] = 14'b11111111111111;

	assign font[0][194] = 14'b11111111111111;
	assign font[1][194] = 14'b11111111111111;
	assign font[2][194] = 14'b11111111111111;
	assign font[3][194] = 14'b11111111111111;
	assign font[4][194] = 14'b11111111111111;
	assign font[5][194] = 14'b11111111111111;
	assign font[6][194] = 14'b11111111111111;
	assign font[7][194] = 14'b11111111111111;
	assign font[8][194] = 14'b11111111111111;
	assign font[9][194] = 14'b11111111111111;
	assign font[10][194] = 14'b11111111111111;
	assign font[11][194] = 14'b11111111111111;
	assign font[12][194] = 14'b11111111111111;
	assign font[13][194] = 14'b11111111111111;
	assign font[14][194] = 14'b11111111111111;
	assign font[15][194] = 14'b11111111111111;
	assign font[16][194] = 14'b11111111111111;
	assign font[17][194] = 14'b11111111111111;
	assign font[18][194] = 14'b11111111111111;
	assign font[19][194] = 14'b11111111111111;
	assign font[20][194] = 14'b11111111111111;
	assign font[21][194] = 14'b11111111111111;
	assign font[22][194] = 14'b11111111111111;
	assign font[23][194] = 14'b11111111111111;
	assign font[24][194] = 14'b11111111111111;
	assign font[25][194] = 14'b11111111111111;
	assign font[26][194] = 14'b11111111111111;
	assign font[27][194] = 14'b11111111111111;
	assign font[28][194] = 14'b11111111111111;
	assign font[29][194] = 14'b11111111111111;
	assign font[30][194] = 14'b11111111111111;
	assign font[31][194] = 14'b11111111111111;

	assign font[0][195] = 14'b11111111111111;
	assign font[1][195] = 14'b11111111111111;
	assign font[2][195] = 14'b11111111111111;
	assign font[3][195] = 14'b11111111111111;
	assign font[4][195] = 14'b11111111111111;
	assign font[5][195] = 14'b11111111111111;
	assign font[6][195] = 14'b11111111111111;
	assign font[7][195] = 14'b11111111111111;
	assign font[8][195] = 14'b11111111111111;
	assign font[9][195] = 14'b11111111111111;
	assign font[10][195] = 14'b11111111111111;
	assign font[11][195] = 14'b11111111111111;
	assign font[12][195] = 14'b11111111111111;
	assign font[13][195] = 14'b11111111111111;
	assign font[14][195] = 14'b11111111111111;
	assign font[15][195] = 14'b11111111111111;
	assign font[16][195] = 14'b11111111111111;
	assign font[17][195] = 14'b11111111111111;
	assign font[18][195] = 14'b11111111111111;
	assign font[19][195] = 14'b11111111111111;
	assign font[20][195] = 14'b11111111111111;
	assign font[21][195] = 14'b11111111111111;
	assign font[22][195] = 14'b11111111111111;
	assign font[23][195] = 14'b11111111111111;
	assign font[24][195] = 14'b11111111111111;
	assign font[25][195] = 14'b11111111111111;
	assign font[26][195] = 14'b11111111111111;
	assign font[27][195] = 14'b11111111111111;
	assign font[28][195] = 14'b11111111111111;
	assign font[29][195] = 14'b11111111111111;
	assign font[30][195] = 14'b11111111111111;
	assign font[31][195] = 14'b11111111111111;

	assign font[0][196] = 14'b11111111111111;
	assign font[1][196] = 14'b11111111111111;
	assign font[2][196] = 14'b11111111111111;
	assign font[3][196] = 14'b11111111111111;
	assign font[4][196] = 14'b11111111111111;
	assign font[5][196] = 14'b11111111111111;
	assign font[6][196] = 14'b11111111111111;
	assign font[7][196] = 14'b11111111111111;
	assign font[8][196] = 14'b11111111111111;
	assign font[9][196] = 14'b11111111111111;
	assign font[10][196] = 14'b11111111111111;
	assign font[11][196] = 14'b11111111111111;
	assign font[12][196] = 14'b11111111111111;
	assign font[13][196] = 14'b11111111111111;
	assign font[14][196] = 14'b11111111111111;
	assign font[15][196] = 14'b11111111111111;
	assign font[16][196] = 14'b11111111111111;
	assign font[17][196] = 14'b11111111111111;
	assign font[18][196] = 14'b11111111111111;
	assign font[19][196] = 14'b11111111111111;
	assign font[20][196] = 14'b11111111111111;
	assign font[21][196] = 14'b11111111111111;
	assign font[22][196] = 14'b11111111111111;
	assign font[23][196] = 14'b11111111111111;
	assign font[24][196] = 14'b11111111111111;
	assign font[25][196] = 14'b11111111111111;
	assign font[26][196] = 14'b11111111111111;
	assign font[27][196] = 14'b11111111111111;
	assign font[28][196] = 14'b11111111111111;
	assign font[29][196] = 14'b11111111111111;
	assign font[30][196] = 14'b11111111111111;
	assign font[31][196] = 14'b11111111111111;

	assign font[0][197] = 14'b11111111111111;
	assign font[1][197] = 14'b11111111111111;
	assign font[2][197] = 14'b11111111111111;
	assign font[3][197] = 14'b11111111111111;
	assign font[4][197] = 14'b11111111111111;
	assign font[5][197] = 14'b11111111111111;
	assign font[6][197] = 14'b11111111111111;
	assign font[7][197] = 14'b11111111111111;
	assign font[8][197] = 14'b11111111111111;
	assign font[9][197] = 14'b11111111111111;
	assign font[10][197] = 14'b11111111111111;
	assign font[11][197] = 14'b11111111111111;
	assign font[12][197] = 14'b11111111111111;
	assign font[13][197] = 14'b11111111111111;
	assign font[14][197] = 14'b11111111111111;
	assign font[15][197] = 14'b11111111111111;
	assign font[16][197] = 14'b11111111111111;
	assign font[17][197] = 14'b11111111111111;
	assign font[18][197] = 14'b11111111111111;
	assign font[19][197] = 14'b11111111111111;
	assign font[20][197] = 14'b11111111111111;
	assign font[21][197] = 14'b11111111111111;
	assign font[22][197] = 14'b11111111111111;
	assign font[23][197] = 14'b11111111111111;
	assign font[24][197] = 14'b11111111111111;
	assign font[25][197] = 14'b11111111111111;
	assign font[26][197] = 14'b11111111111111;
	assign font[27][197] = 14'b11111111111111;
	assign font[28][197] = 14'b11111111111111;
	assign font[29][197] = 14'b11111111111111;
	assign font[30][197] = 14'b11111111111111;
	assign font[31][197] = 14'b11111111111111;

	assign font[0][198] = 14'b11111111111111;
	assign font[1][198] = 14'b11111111111111;
	assign font[2][198] = 14'b11111111111111;
	assign font[3][198] = 14'b11111111111111;
	assign font[4][198] = 14'b11111111111111;
	assign font[5][198] = 14'b11111111111111;
	assign font[6][198] = 14'b11111111111111;
	assign font[7][198] = 14'b11111111111111;
	assign font[8][198] = 14'b11111111111111;
	assign font[9][198] = 14'b11111111111111;
	assign font[10][198] = 14'b11111111111111;
	assign font[11][198] = 14'b11111111111111;
	assign font[12][198] = 14'b11111111111111;
	assign font[13][198] = 14'b11111111111111;
	assign font[14][198] = 14'b11111111111111;
	assign font[15][198] = 14'b11111111111111;
	assign font[16][198] = 14'b11111111111111;
	assign font[17][198] = 14'b11111111111111;
	assign font[18][198] = 14'b11111111111111;
	assign font[19][198] = 14'b11111111111111;
	assign font[20][198] = 14'b11111111111111;
	assign font[21][198] = 14'b11111111111111;
	assign font[22][198] = 14'b11111111111111;
	assign font[23][198] = 14'b11111111111111;
	assign font[24][198] = 14'b11111111111111;
	assign font[25][198] = 14'b11111111111111;
	assign font[26][198] = 14'b11111111111111;
	assign font[27][198] = 14'b11111111111111;
	assign font[28][198] = 14'b11111111111111;
	assign font[29][198] = 14'b11111111111111;
	assign font[30][198] = 14'b11111111111111;
	assign font[31][198] = 14'b11111111111111;

	assign font[0][199] = 14'b11111111111111;
	assign font[1][199] = 14'b11111111111111;
	assign font[2][199] = 14'b11111111111111;
	assign font[3][199] = 14'b11111111111111;
	assign font[4][199] = 14'b11111111111111;
	assign font[5][199] = 14'b11111111111111;
	assign font[6][199] = 14'b11111111111111;
	assign font[7][199] = 14'b11111111111111;
	assign font[8][199] = 14'b11111111111111;
	assign font[9][199] = 14'b11111111111111;
	assign font[10][199] = 14'b11111111111111;
	assign font[11][199] = 14'b11111111111111;
	assign font[12][199] = 14'b11111111111111;
	assign font[13][199] = 14'b11111111111111;
	assign font[14][199] = 14'b11111111111111;
	assign font[15][199] = 14'b11111111111111;
	assign font[16][199] = 14'b11111111111111;
	assign font[17][199] = 14'b11111111111111;
	assign font[18][199] = 14'b11111111111111;
	assign font[19][199] = 14'b11111111111111;
	assign font[20][199] = 14'b11111111111111;
	assign font[21][199] = 14'b11111111111111;
	assign font[22][199] = 14'b11111111111111;
	assign font[23][199] = 14'b11111111111111;
	assign font[24][199] = 14'b11111111111111;
	assign font[25][199] = 14'b11111111111111;
	assign font[26][199] = 14'b11111111111111;
	assign font[27][199] = 14'b11111111111111;
	assign font[28][199] = 14'b11111111111111;
	assign font[29][199] = 14'b11111111111111;
	assign font[30][199] = 14'b11111111111111;
	assign font[31][199] = 14'b11111111111111;

	assign font[0][200] = 14'b11111111111111;
	assign font[1][200] = 14'b11111111111111;
	assign font[2][200] = 14'b11111111111111;
	assign font[3][200] = 14'b11111111111111;
	assign font[4][200] = 14'b11111111111111;
	assign font[5][200] = 14'b11111111111111;
	assign font[6][200] = 14'b11111111111111;
	assign font[7][200] = 14'b11111111111111;
	assign font[8][200] = 14'b11111111111111;
	assign font[9][200] = 14'b11111111111111;
	assign font[10][200] = 14'b11111111111111;
	assign font[11][200] = 14'b11111111111111;
	assign font[12][200] = 14'b11111111111111;
	assign font[13][200] = 14'b11111111111111;
	assign font[14][200] = 14'b11111111111111;
	assign font[15][200] = 14'b11111111111111;
	assign font[16][200] = 14'b11111111111111;
	assign font[17][200] = 14'b11111111111111;
	assign font[18][200] = 14'b11111111111111;
	assign font[19][200] = 14'b11111111111111;
	assign font[20][200] = 14'b11111111111111;
	assign font[21][200] = 14'b11111111111111;
	assign font[22][200] = 14'b11111111111111;
	assign font[23][200] = 14'b11111111111111;
	assign font[24][200] = 14'b11111111111111;
	assign font[25][200] = 14'b11111111111111;
	assign font[26][200] = 14'b11111111111111;
	assign font[27][200] = 14'b11111111111111;
	assign font[28][200] = 14'b11111111111111;
	assign font[29][200] = 14'b11111111111111;
	assign font[30][200] = 14'b11111111111111;
	assign font[31][200] = 14'b11111111111111;

	assign font[0][201] = 14'b11111111111111;
	assign font[1][201] = 14'b11111111111111;
	assign font[2][201] = 14'b11111111111111;
	assign font[3][201] = 14'b11111111111111;
	assign font[4][201] = 14'b11111111111111;
	assign font[5][201] = 14'b11111111111111;
	assign font[6][201] = 14'b11111111111111;
	assign font[7][201] = 14'b11111111111111;
	assign font[8][201] = 14'b11111111111111;
	assign font[9][201] = 14'b11111111111111;
	assign font[10][201] = 14'b11111111111111;
	assign font[11][201] = 14'b11111111111111;
	assign font[12][201] = 14'b11111111111111;
	assign font[13][201] = 14'b11111111111111;
	assign font[14][201] = 14'b11111111111111;
	assign font[15][201] = 14'b11111111111111;
	assign font[16][201] = 14'b11111111111111;
	assign font[17][201] = 14'b11111111111111;
	assign font[18][201] = 14'b11111111111111;
	assign font[19][201] = 14'b11111111111111;
	assign font[20][201] = 14'b11111111111111;
	assign font[21][201] = 14'b11111111111111;
	assign font[22][201] = 14'b11111111111111;
	assign font[23][201] = 14'b11111111111111;
	assign font[24][201] = 14'b11111111111111;
	assign font[25][201] = 14'b11111111111111;
	assign font[26][201] = 14'b11111111111111;
	assign font[27][201] = 14'b11111111111111;
	assign font[28][201] = 14'b11111111111111;
	assign font[29][201] = 14'b11111111111111;
	assign font[30][201] = 14'b11111111111111;
	assign font[31][201] = 14'b11111111111111;

	assign font[0][202] = 14'b11111111111111;
	assign font[1][202] = 14'b11111111111111;
	assign font[2][202] = 14'b11111111111111;
	assign font[3][202] = 14'b11111111111111;
	assign font[4][202] = 14'b11111111111111;
	assign font[5][202] = 14'b11111111111111;
	assign font[6][202] = 14'b11111111111111;
	assign font[7][202] = 14'b11111111111111;
	assign font[8][202] = 14'b11111111111111;
	assign font[9][202] = 14'b11111111111111;
	assign font[10][202] = 14'b11111111111111;
	assign font[11][202] = 14'b11111111111111;
	assign font[12][202] = 14'b11111111111111;
	assign font[13][202] = 14'b11111111111111;
	assign font[14][202] = 14'b11111111111111;
	assign font[15][202] = 14'b11111111111111;
	assign font[16][202] = 14'b11111111111111;
	assign font[17][202] = 14'b11111111111111;
	assign font[18][202] = 14'b11111111111111;
	assign font[19][202] = 14'b11111111111111;
	assign font[20][202] = 14'b11111111111111;
	assign font[21][202] = 14'b11111111111111;
	assign font[22][202] = 14'b11111111111111;
	assign font[23][202] = 14'b11111111111111;
	assign font[24][202] = 14'b11111111111111;
	assign font[25][202] = 14'b11111111111111;
	assign font[26][202] = 14'b11111111111111;
	assign font[27][202] = 14'b11111111111111;
	assign font[28][202] = 14'b11111111111111;
	assign font[29][202] = 14'b11111111111111;
	assign font[30][202] = 14'b11111111111111;
	assign font[31][202] = 14'b11111111111111;

	assign font[0][203] = 14'b11111111111111;
	assign font[1][203] = 14'b11111111111111;
	assign font[2][203] = 14'b11111111111111;
	assign font[3][203] = 14'b11111111111111;
	assign font[4][203] = 14'b11111111111111;
	assign font[5][203] = 14'b11111111111111;
	assign font[6][203] = 14'b11111111111111;
	assign font[7][203] = 14'b11111111111111;
	assign font[8][203] = 14'b11111111111111;
	assign font[9][203] = 14'b11111111111111;
	assign font[10][203] = 14'b11111111111111;
	assign font[11][203] = 14'b11111111111111;
	assign font[12][203] = 14'b11111111111111;
	assign font[13][203] = 14'b11111111111111;
	assign font[14][203] = 14'b11111111111111;
	assign font[15][203] = 14'b11111111111111;
	assign font[16][203] = 14'b11111111111111;
	assign font[17][203] = 14'b11111111111111;
	assign font[18][203] = 14'b11111111111111;
	assign font[19][203] = 14'b11111111111111;
	assign font[20][203] = 14'b11111111111111;
	assign font[21][203] = 14'b11111111111111;
	assign font[22][203] = 14'b11111111111111;
	assign font[23][203] = 14'b11111111111111;
	assign font[24][203] = 14'b11111111111111;
	assign font[25][203] = 14'b11111111111111;
	assign font[26][203] = 14'b11111111111111;
	assign font[27][203] = 14'b11111111111111;
	assign font[28][203] = 14'b11111111111111;
	assign font[29][203] = 14'b11111111111111;
	assign font[30][203] = 14'b11111111111111;
	assign font[31][203] = 14'b11111111111111;

	assign font[0][204] = 14'b11111111111111;
	assign font[1][204] = 14'b11111111111111;
	assign font[2][204] = 14'b11111111111111;
	assign font[3][204] = 14'b11111111111111;
	assign font[4][204] = 14'b11111111111111;
	assign font[5][204] = 14'b11111111111111;
	assign font[6][204] = 14'b11111111111111;
	assign font[7][204] = 14'b11111111111111;
	assign font[8][204] = 14'b11111111111111;
	assign font[9][204] = 14'b11111111111111;
	assign font[10][204] = 14'b11111111111111;
	assign font[11][204] = 14'b11111111111111;
	assign font[12][204] = 14'b11111111111111;
	assign font[13][204] = 14'b11111111111111;
	assign font[14][204] = 14'b11111111111111;
	assign font[15][204] = 14'b11111111111111;
	assign font[16][204] = 14'b11111111111111;
	assign font[17][204] = 14'b11111111111111;
	assign font[18][204] = 14'b11111111111111;
	assign font[19][204] = 14'b11111111111111;
	assign font[20][204] = 14'b11111111111111;
	assign font[21][204] = 14'b11111111111111;
	assign font[22][204] = 14'b11111111111111;
	assign font[23][204] = 14'b11111111111111;
	assign font[24][204] = 14'b11111111111111;
	assign font[25][204] = 14'b11111111111111;
	assign font[26][204] = 14'b11111111111111;
	assign font[27][204] = 14'b11111111111111;
	assign font[28][204] = 14'b11111111111111;
	assign font[29][204] = 14'b11111111111111;
	assign font[30][204] = 14'b11111111111111;
	assign font[31][204] = 14'b11111111111111;

	assign font[0][205] = 14'b11111111111111;
	assign font[1][205] = 14'b11111111111111;
	assign font[2][205] = 14'b11111111111111;
	assign font[3][205] = 14'b11111111111111;
	assign font[4][205] = 14'b11111111111111;
	assign font[5][205] = 14'b11111111111111;
	assign font[6][205] = 14'b11111111111111;
	assign font[7][205] = 14'b11111111111111;
	assign font[8][205] = 14'b11111111111111;
	assign font[9][205] = 14'b11111111111111;
	assign font[10][205] = 14'b11111111111111;
	assign font[11][205] = 14'b11111111111111;
	assign font[12][205] = 14'b11111111111111;
	assign font[13][205] = 14'b11111111111111;
	assign font[14][205] = 14'b11111111111111;
	assign font[15][205] = 14'b11111111111111;
	assign font[16][205] = 14'b11111111111111;
	assign font[17][205] = 14'b11111111111111;
	assign font[18][205] = 14'b11111111111111;
	assign font[19][205] = 14'b11111111111111;
	assign font[20][205] = 14'b11111111111111;
	assign font[21][205] = 14'b11111111111111;
	assign font[22][205] = 14'b11111111111111;
	assign font[23][205] = 14'b11111111111111;
	assign font[24][205] = 14'b11111111111111;
	assign font[25][205] = 14'b11111111111111;
	assign font[26][205] = 14'b11111111111111;
	assign font[27][205] = 14'b11111111111111;
	assign font[28][205] = 14'b11111111111111;
	assign font[29][205] = 14'b11111111111111;
	assign font[30][205] = 14'b11111111111111;
	assign font[31][205] = 14'b11111111111111;

	assign font[0][206] = 14'b11111111111111;
	assign font[1][206] = 14'b11111111111111;
	assign font[2][206] = 14'b11111111111111;
	assign font[3][206] = 14'b11111111111111;
	assign font[4][206] = 14'b11111111111111;
	assign font[5][206] = 14'b11111111111111;
	assign font[6][206] = 14'b11111111111111;
	assign font[7][206] = 14'b11111111111111;
	assign font[8][206] = 14'b11111111111111;
	assign font[9][206] = 14'b11111111111111;
	assign font[10][206] = 14'b11111111111111;
	assign font[11][206] = 14'b11111111111111;
	assign font[12][206] = 14'b11111111111111;
	assign font[13][206] = 14'b11111111111111;
	assign font[14][206] = 14'b11111111111111;
	assign font[15][206] = 14'b11111111111111;
	assign font[16][206] = 14'b11111111111111;
	assign font[17][206] = 14'b11111111111111;
	assign font[18][206] = 14'b11111111111111;
	assign font[19][206] = 14'b11111111111111;
	assign font[20][206] = 14'b11111111111111;
	assign font[21][206] = 14'b11111111111111;
	assign font[22][206] = 14'b11111111111111;
	assign font[23][206] = 14'b11111111111111;
	assign font[24][206] = 14'b11111111111111;
	assign font[25][206] = 14'b11111111111111;
	assign font[26][206] = 14'b11111111111111;
	assign font[27][206] = 14'b11111111111111;
	assign font[28][206] = 14'b11111111111111;
	assign font[29][206] = 14'b11111111111111;
	assign font[30][206] = 14'b11111111111111;
	assign font[31][206] = 14'b11111111111111;

	assign font[0][207] = 14'b11111111111111;
	assign font[1][207] = 14'b11111111111111;
	assign font[2][207] = 14'b11111111111111;
	assign font[3][207] = 14'b11111111111111;
	assign font[4][207] = 14'b11111111111111;
	assign font[5][207] = 14'b11111111111111;
	assign font[6][207] = 14'b11111111111111;
	assign font[7][207] = 14'b11111111111111;
	assign font[8][207] = 14'b11111111111111;
	assign font[9][207] = 14'b11111111111111;
	assign font[10][207] = 14'b11111111111111;
	assign font[11][207] = 14'b11111111111111;
	assign font[12][207] = 14'b11111111111111;
	assign font[13][207] = 14'b11111111111111;
	assign font[14][207] = 14'b11111111111111;
	assign font[15][207] = 14'b11111111111111;
	assign font[16][207] = 14'b11111111111111;
	assign font[17][207] = 14'b11111111111111;
	assign font[18][207] = 14'b11111111111111;
	assign font[19][207] = 14'b11111111111111;
	assign font[20][207] = 14'b11111111111111;
	assign font[21][207] = 14'b11111111111111;
	assign font[22][207] = 14'b11111111111111;
	assign font[23][207] = 14'b11111111111111;
	assign font[24][207] = 14'b11111111111111;
	assign font[25][207] = 14'b11111111111111;
	assign font[26][207] = 14'b11111111111111;
	assign font[27][207] = 14'b11111111111111;
	assign font[28][207] = 14'b11111111111111;
	assign font[29][207] = 14'b11111111111111;
	assign font[30][207] = 14'b11111111111111;
	assign font[31][207] = 14'b11111111111111;

	assign font[0][208] = 14'b11111111111111;
	assign font[1][208] = 14'b11111111111111;
	assign font[2][208] = 14'b11111111111111;
	assign font[3][208] = 14'b11111111111111;
	assign font[4][208] = 14'b11111111111111;
	assign font[5][208] = 14'b11111111111111;
	assign font[6][208] = 14'b11111111111111;
	assign font[7][208] = 14'b11111111111111;
	assign font[8][208] = 14'b11111111111111;
	assign font[9][208] = 14'b11111111111111;
	assign font[10][208] = 14'b11111111111111;
	assign font[11][208] = 14'b11111111111111;
	assign font[12][208] = 14'b11111111111111;
	assign font[13][208] = 14'b11111111111111;
	assign font[14][208] = 14'b11111111111111;
	assign font[15][208] = 14'b11111111111111;
	assign font[16][208] = 14'b11111111111111;
	assign font[17][208] = 14'b11111111111111;
	assign font[18][208] = 14'b11111111111111;
	assign font[19][208] = 14'b11111111111111;
	assign font[20][208] = 14'b11111111111111;
	assign font[21][208] = 14'b11111111111111;
	assign font[22][208] = 14'b11111111111111;
	assign font[23][208] = 14'b11111111111111;
	assign font[24][208] = 14'b11111111111111;
	assign font[25][208] = 14'b11111111111111;
	assign font[26][208] = 14'b11111111111111;
	assign font[27][208] = 14'b11111111111111;
	assign font[28][208] = 14'b11111111111111;
	assign font[29][208] = 14'b11111111111111;
	assign font[30][208] = 14'b11111111111111;
	assign font[31][208] = 14'b11111111111111;

	assign font[0][209] = 14'b11111111111111;
	assign font[1][209] = 14'b11111111111111;
	assign font[2][209] = 14'b11111111111111;
	assign font[3][209] = 14'b11111111111111;
	assign font[4][209] = 14'b11111111111111;
	assign font[5][209] = 14'b11111111111111;
	assign font[6][209] = 14'b11111111111111;
	assign font[7][209] = 14'b11111111111111;
	assign font[8][209] = 14'b11111111111111;
	assign font[9][209] = 14'b11111111111111;
	assign font[10][209] = 14'b11111111111111;
	assign font[11][209] = 14'b11111111111111;
	assign font[12][209] = 14'b11111111111111;
	assign font[13][209] = 14'b11111111111111;
	assign font[14][209] = 14'b11111111111111;
	assign font[15][209] = 14'b11111111111111;
	assign font[16][209] = 14'b11111111111111;
	assign font[17][209] = 14'b11111111111111;
	assign font[18][209] = 14'b11111111111111;
	assign font[19][209] = 14'b11111111111111;
	assign font[20][209] = 14'b11111111111111;
	assign font[21][209] = 14'b11111111111111;
	assign font[22][209] = 14'b11111111111111;
	assign font[23][209] = 14'b11111111111111;
	assign font[24][209] = 14'b11111111111111;
	assign font[25][209] = 14'b11111111111111;
	assign font[26][209] = 14'b11111111111111;
	assign font[27][209] = 14'b11111111111111;
	assign font[28][209] = 14'b11111111111111;
	assign font[29][209] = 14'b11111111111111;
	assign font[30][209] = 14'b11111111111111;
	assign font[31][209] = 14'b11111111111111;

	assign font[0][210] = 14'b11111111111111;
	assign font[1][210] = 14'b11111111111111;
	assign font[2][210] = 14'b11111111111111;
	assign font[3][210] = 14'b11111111111111;
	assign font[4][210] = 14'b11111111111111;
	assign font[5][210] = 14'b11111111111111;
	assign font[6][210] = 14'b11111111111111;
	assign font[7][210] = 14'b11111111111111;
	assign font[8][210] = 14'b11111111111111;
	assign font[9][210] = 14'b11111111111111;
	assign font[10][210] = 14'b11111111111111;
	assign font[11][210] = 14'b11111111111111;
	assign font[12][210] = 14'b11111111111111;
	assign font[13][210] = 14'b11111111111111;
	assign font[14][210] = 14'b11111111111111;
	assign font[15][210] = 14'b11111111111111;
	assign font[16][210] = 14'b11111111111111;
	assign font[17][210] = 14'b11111111111111;
	assign font[18][210] = 14'b11111111111111;
	assign font[19][210] = 14'b11111111111111;
	assign font[20][210] = 14'b11111111111111;
	assign font[21][210] = 14'b11111111111111;
	assign font[22][210] = 14'b11111111111111;
	assign font[23][210] = 14'b11111111111111;
	assign font[24][210] = 14'b11111111111111;
	assign font[25][210] = 14'b11111111111111;
	assign font[26][210] = 14'b11111111111111;
	assign font[27][210] = 14'b11111111111111;
	assign font[28][210] = 14'b11111111111111;
	assign font[29][210] = 14'b11111111111111;
	assign font[30][210] = 14'b11111111111111;
	assign font[31][210] = 14'b11111111111111;

	assign font[0][211] = 14'b11111111111111;
	assign font[1][211] = 14'b11111111111111;
	assign font[2][211] = 14'b11111111111111;
	assign font[3][211] = 14'b11111111111111;
	assign font[4][211] = 14'b11111111111111;
	assign font[5][211] = 14'b11111111111111;
	assign font[6][211] = 14'b11111111111111;
	assign font[7][211] = 14'b11111111111111;
	assign font[8][211] = 14'b11111111111111;
	assign font[9][211] = 14'b11111111111111;
	assign font[10][211] = 14'b11111111111111;
	assign font[11][211] = 14'b11111111111111;
	assign font[12][211] = 14'b11111111111111;
	assign font[13][211] = 14'b11111111111111;
	assign font[14][211] = 14'b11111111111111;
	assign font[15][211] = 14'b11111111111111;
	assign font[16][211] = 14'b11111111111111;
	assign font[17][211] = 14'b11111111111111;
	assign font[18][211] = 14'b11111111111111;
	assign font[19][211] = 14'b11111111111111;
	assign font[20][211] = 14'b11111111111111;
	assign font[21][211] = 14'b11111111111111;
	assign font[22][211] = 14'b11111111111111;
	assign font[23][211] = 14'b11111111111111;
	assign font[24][211] = 14'b11111111111111;
	assign font[25][211] = 14'b11111111111111;
	assign font[26][211] = 14'b11111111111111;
	assign font[27][211] = 14'b11111111111111;
	assign font[28][211] = 14'b11111111111111;
	assign font[29][211] = 14'b11111111111111;
	assign font[30][211] = 14'b11111111111111;
	assign font[31][211] = 14'b11111111111111;

	assign font[0][212] = 14'b11111111111111;
	assign font[1][212] = 14'b11111111111111;
	assign font[2][212] = 14'b11111111111111;
	assign font[3][212] = 14'b11111111111111;
	assign font[4][212] = 14'b11111111111111;
	assign font[5][212] = 14'b11111111111111;
	assign font[6][212] = 14'b11111111111111;
	assign font[7][212] = 14'b11111111111111;
	assign font[8][212] = 14'b11111111111111;
	assign font[9][212] = 14'b11111111111111;
	assign font[10][212] = 14'b11111111111111;
	assign font[11][212] = 14'b11111111111111;
	assign font[12][212] = 14'b11111111111111;
	assign font[13][212] = 14'b11111111111111;
	assign font[14][212] = 14'b11111111111111;
	assign font[15][212] = 14'b11111111111111;
	assign font[16][212] = 14'b11111111111111;
	assign font[17][212] = 14'b11111111111111;
	assign font[18][212] = 14'b11111111111111;
	assign font[19][212] = 14'b11111111111111;
	assign font[20][212] = 14'b11111111111111;
	assign font[21][212] = 14'b11111111111111;
	assign font[22][212] = 14'b11111111111111;
	assign font[23][212] = 14'b11111111111111;
	assign font[24][212] = 14'b11111111111111;
	assign font[25][212] = 14'b11111111111111;
	assign font[26][212] = 14'b11111111111111;
	assign font[27][212] = 14'b11111111111111;
	assign font[28][212] = 14'b11111111111111;
	assign font[29][212] = 14'b11111111111111;
	assign font[30][212] = 14'b11111111111111;
	assign font[31][212] = 14'b11111111111111;

	assign font[0][213] = 14'b11111111111111;
	assign font[1][213] = 14'b11111111111111;
	assign font[2][213] = 14'b11111111111111;
	assign font[3][213] = 14'b11111111111111;
	assign font[4][213] = 14'b11111111111111;
	assign font[5][213] = 14'b11111111111111;
	assign font[6][213] = 14'b11111111111111;
	assign font[7][213] = 14'b11111111111111;
	assign font[8][213] = 14'b11111111111111;
	assign font[9][213] = 14'b11111111111111;
	assign font[10][213] = 14'b11111111111111;
	assign font[11][213] = 14'b11111111111111;
	assign font[12][213] = 14'b11111111111111;
	assign font[13][213] = 14'b11111111111111;
	assign font[14][213] = 14'b11111111111111;
	assign font[15][213] = 14'b11111111111111;
	assign font[16][213] = 14'b11111111111111;
	assign font[17][213] = 14'b11111111111111;
	assign font[18][213] = 14'b11111111111111;
	assign font[19][213] = 14'b11111111111111;
	assign font[20][213] = 14'b11111111111111;
	assign font[21][213] = 14'b11111111111111;
	assign font[22][213] = 14'b11111111111111;
	assign font[23][213] = 14'b11111111111111;
	assign font[24][213] = 14'b11111111111111;
	assign font[25][213] = 14'b11111111111111;
	assign font[26][213] = 14'b11111111111111;
	assign font[27][213] = 14'b11111111111111;
	assign font[28][213] = 14'b11111111111111;
	assign font[29][213] = 14'b11111111111111;
	assign font[30][213] = 14'b11111111111111;
	assign font[31][213] = 14'b11111111111111;

	assign font[0][214] = 14'b11111111111111;
	assign font[1][214] = 14'b11111111111111;
	assign font[2][214] = 14'b11111111111111;
	assign font[3][214] = 14'b11111111111111;
	assign font[4][214] = 14'b11111111111111;
	assign font[5][214] = 14'b11111111111111;
	assign font[6][214] = 14'b11111111111111;
	assign font[7][214] = 14'b11111111111111;
	assign font[8][214] = 14'b11111111111111;
	assign font[9][214] = 14'b11111111111111;
	assign font[10][214] = 14'b11111111111111;
	assign font[11][214] = 14'b11111111111111;
	assign font[12][214] = 14'b11111111111111;
	assign font[13][214] = 14'b11111111111111;
	assign font[14][214] = 14'b11111111111111;
	assign font[15][214] = 14'b11111111111111;
	assign font[16][214] = 14'b11111111111111;
	assign font[17][214] = 14'b11111111111111;
	assign font[18][214] = 14'b11111111111111;
	assign font[19][214] = 14'b11111111111111;
	assign font[20][214] = 14'b11111111111111;
	assign font[21][214] = 14'b11111111111111;
	assign font[22][214] = 14'b11111111111111;
	assign font[23][214] = 14'b11111111111111;
	assign font[24][214] = 14'b11111111111111;
	assign font[25][214] = 14'b11111111111111;
	assign font[26][214] = 14'b11111111111111;
	assign font[27][214] = 14'b11111111111111;
	assign font[28][214] = 14'b11111111111111;
	assign font[29][214] = 14'b11111111111111;
	assign font[30][214] = 14'b11111111111111;
	assign font[31][214] = 14'b11111111111111;

	assign font[0][215] = 14'b11111111111111;
	assign font[1][215] = 14'b11111111111111;
	assign font[2][215] = 14'b11111111111111;
	assign font[3][215] = 14'b11111111111111;
	assign font[4][215] = 14'b11111111111111;
	assign font[5][215] = 14'b11111111111111;
	assign font[6][215] = 14'b11111111111111;
	assign font[7][215] = 14'b11111111111111;
	assign font[8][215] = 14'b11111111111111;
	assign font[9][215] = 14'b11111111111111;
	assign font[10][215] = 14'b11111111111111;
	assign font[11][215] = 14'b11111111111111;
	assign font[12][215] = 14'b11111111111111;
	assign font[13][215] = 14'b11111111111111;
	assign font[14][215] = 14'b11111111111111;
	assign font[15][215] = 14'b11111111111111;
	assign font[16][215] = 14'b11111111111111;
	assign font[17][215] = 14'b11111111111111;
	assign font[18][215] = 14'b11111111111111;
	assign font[19][215] = 14'b11111111111111;
	assign font[20][215] = 14'b11111111111111;
	assign font[21][215] = 14'b11111111111111;
	assign font[22][215] = 14'b11111111111111;
	assign font[23][215] = 14'b11111111111111;
	assign font[24][215] = 14'b11111111111111;
	assign font[25][215] = 14'b11111111111111;
	assign font[26][215] = 14'b11111111111111;
	assign font[27][215] = 14'b11111111111111;
	assign font[28][215] = 14'b11111111111111;
	assign font[29][215] = 14'b11111111111111;
	assign font[30][215] = 14'b11111111111111;
	assign font[31][215] = 14'b11111111111111;

	assign font[0][216] = 14'b11111111111111;
	assign font[1][216] = 14'b11111111111111;
	assign font[2][216] = 14'b11111111111111;
	assign font[3][216] = 14'b11111111111111;
	assign font[4][216] = 14'b11111111111111;
	assign font[5][216] = 14'b11111111111111;
	assign font[6][216] = 14'b11111111111111;
	assign font[7][216] = 14'b11111111111111;
	assign font[8][216] = 14'b11111111111111;
	assign font[9][216] = 14'b11111111111111;
	assign font[10][216] = 14'b11111111111111;
	assign font[11][216] = 14'b11111111111111;
	assign font[12][216] = 14'b11111111111111;
	assign font[13][216] = 14'b11111111111111;
	assign font[14][216] = 14'b11111111111111;
	assign font[15][216] = 14'b11111111111111;
	assign font[16][216] = 14'b11111111111111;
	assign font[17][216] = 14'b11111111111111;
	assign font[18][216] = 14'b11111111111111;
	assign font[19][216] = 14'b11111111111111;
	assign font[20][216] = 14'b11111111111111;
	assign font[21][216] = 14'b11111111111111;
	assign font[22][216] = 14'b11111111111111;
	assign font[23][216] = 14'b11111111111111;
	assign font[24][216] = 14'b11111111111111;
	assign font[25][216] = 14'b11111111111111;
	assign font[26][216] = 14'b11111111111111;
	assign font[27][216] = 14'b11111111111111;
	assign font[28][216] = 14'b11111111111111;
	assign font[29][216] = 14'b11111111111111;
	assign font[30][216] = 14'b11111111111111;
	assign font[31][216] = 14'b11111111111111;

	assign font[0][217] = 14'b11111111111111;
	assign font[1][217] = 14'b11111111111111;
	assign font[2][217] = 14'b11111111111111;
	assign font[3][217] = 14'b11111111111111;
	assign font[4][217] = 14'b11111111111111;
	assign font[5][217] = 14'b11111111111111;
	assign font[6][217] = 14'b11111111111111;
	assign font[7][217] = 14'b11111111111111;
	assign font[8][217] = 14'b11111111111111;
	assign font[9][217] = 14'b11111111111111;
	assign font[10][217] = 14'b11111111111111;
	assign font[11][217] = 14'b11111111111111;
	assign font[12][217] = 14'b11111111111111;
	assign font[13][217] = 14'b11111111111111;
	assign font[14][217] = 14'b11111111111111;
	assign font[15][217] = 14'b11111111111111;
	assign font[16][217] = 14'b11111111111111;
	assign font[17][217] = 14'b11111111111111;
	assign font[18][217] = 14'b11111111111111;
	assign font[19][217] = 14'b11111111111111;
	assign font[20][217] = 14'b11111111111111;
	assign font[21][217] = 14'b11111111111111;
	assign font[22][217] = 14'b11111111111111;
	assign font[23][217] = 14'b11111111111111;
	assign font[24][217] = 14'b11111111111111;
	assign font[25][217] = 14'b11111111111111;
	assign font[26][217] = 14'b11111111111111;
	assign font[27][217] = 14'b11111111111111;
	assign font[28][217] = 14'b11111111111111;
	assign font[29][217] = 14'b11111111111111;
	assign font[30][217] = 14'b11111111111111;
	assign font[31][217] = 14'b11111111111111;

	assign font[0][218] = 14'b11111111111111;
	assign font[1][218] = 14'b11111111111111;
	assign font[2][218] = 14'b11111111111111;
	assign font[3][218] = 14'b11111111111111;
	assign font[4][218] = 14'b11111111111111;
	assign font[5][218] = 14'b11111111111111;
	assign font[6][218] = 14'b11111111111111;
	assign font[7][218] = 14'b11111111111111;
	assign font[8][218] = 14'b11111111111111;
	assign font[9][218] = 14'b11111111111111;
	assign font[10][218] = 14'b11111111111111;
	assign font[11][218] = 14'b11111111111111;
	assign font[12][218] = 14'b11111111111111;
	assign font[13][218] = 14'b11111111111111;
	assign font[14][218] = 14'b11111111111111;
	assign font[15][218] = 14'b11111111111111;
	assign font[16][218] = 14'b11111111111111;
	assign font[17][218] = 14'b11111111111111;
	assign font[18][218] = 14'b11111111111111;
	assign font[19][218] = 14'b11111111111111;
	assign font[20][218] = 14'b11111111111111;
	assign font[21][218] = 14'b11111111111111;
	assign font[22][218] = 14'b11111111111111;
	assign font[23][218] = 14'b11111111111111;
	assign font[24][218] = 14'b11111111111111;
	assign font[25][218] = 14'b11111111111111;
	assign font[26][218] = 14'b11111111111111;
	assign font[27][218] = 14'b11111111111111;
	assign font[28][218] = 14'b11111111111111;
	assign font[29][218] = 14'b11111111111111;
	assign font[30][218] = 14'b11111111111111;
	assign font[31][218] = 14'b11111111111111;

	assign font[0][219] = 14'b11111111111111;
	assign font[1][219] = 14'b11111111111111;
	assign font[2][219] = 14'b11111111111111;
	assign font[3][219] = 14'b11111111111111;
	assign font[4][219] = 14'b11111111111111;
	assign font[5][219] = 14'b11111111111111;
	assign font[6][219] = 14'b11111111111111;
	assign font[7][219] = 14'b11111111111111;
	assign font[8][219] = 14'b11111111111111;
	assign font[9][219] = 14'b11111111111111;
	assign font[10][219] = 14'b11111111111111;
	assign font[11][219] = 14'b11111111111111;
	assign font[12][219] = 14'b11111111111111;
	assign font[13][219] = 14'b11111111111111;
	assign font[14][219] = 14'b11111111111111;
	assign font[15][219] = 14'b11111111111111;
	assign font[16][219] = 14'b11111111111111;
	assign font[17][219] = 14'b11111111111111;
	assign font[18][219] = 14'b11111111111111;
	assign font[19][219] = 14'b11111111111111;
	assign font[20][219] = 14'b11111111111111;
	assign font[21][219] = 14'b11111111111111;
	assign font[22][219] = 14'b11111111111111;
	assign font[23][219] = 14'b11111111111111;
	assign font[24][219] = 14'b11111111111111;
	assign font[25][219] = 14'b11111111111111;
	assign font[26][219] = 14'b11111111111111;
	assign font[27][219] = 14'b11111111111111;
	assign font[28][219] = 14'b11111111111111;
	assign font[29][219] = 14'b11111111111111;
	assign font[30][219] = 14'b11111111111111;
	assign font[31][219] = 14'b11111111111111;

	assign font[0][220] = 14'b11111111111111;
	assign font[1][220] = 14'b11111111111111;
	assign font[2][220] = 14'b11111111111111;
	assign font[3][220] = 14'b11111111111111;
	assign font[4][220] = 14'b11111111111111;
	assign font[5][220] = 14'b11111111111111;
	assign font[6][220] = 14'b11111111111111;
	assign font[7][220] = 14'b11111111111111;
	assign font[8][220] = 14'b11111111111111;
	assign font[9][220] = 14'b11111111111111;
	assign font[10][220] = 14'b11111111111111;
	assign font[11][220] = 14'b11111111111111;
	assign font[12][220] = 14'b11111111111111;
	assign font[13][220] = 14'b11111111111111;
	assign font[14][220] = 14'b11111111111111;
	assign font[15][220] = 14'b11111111111111;
	assign font[16][220] = 14'b11111111111111;
	assign font[17][220] = 14'b11111111111111;
	assign font[18][220] = 14'b11111111111111;
	assign font[19][220] = 14'b11111111111111;
	assign font[20][220] = 14'b11111111111111;
	assign font[21][220] = 14'b11111111111111;
	assign font[22][220] = 14'b11111111111111;
	assign font[23][220] = 14'b11111111111111;
	assign font[24][220] = 14'b11111111111111;
	assign font[25][220] = 14'b11111111111111;
	assign font[26][220] = 14'b11111111111111;
	assign font[27][220] = 14'b11111111111111;
	assign font[28][220] = 14'b11111111111111;
	assign font[29][220] = 14'b11111111111111;
	assign font[30][220] = 14'b11111111111111;
	assign font[31][220] = 14'b11111111111111;

	assign font[0][221] = 14'b11111111111111;
	assign font[1][221] = 14'b11111111111111;
	assign font[2][221] = 14'b11111111111111;
	assign font[3][221] = 14'b11111111111111;
	assign font[4][221] = 14'b11111111111111;
	assign font[5][221] = 14'b11111111111111;
	assign font[6][221] = 14'b11111111111111;
	assign font[7][221] = 14'b11111111111111;
	assign font[8][221] = 14'b11111111111111;
	assign font[9][221] = 14'b11111111111111;
	assign font[10][221] = 14'b11111111111111;
	assign font[11][221] = 14'b11111111111111;
	assign font[12][221] = 14'b11111111111111;
	assign font[13][221] = 14'b11111111111111;
	assign font[14][221] = 14'b11111111111111;
	assign font[15][221] = 14'b11111111111111;
	assign font[16][221] = 14'b11111111111111;
	assign font[17][221] = 14'b11111111111111;
	assign font[18][221] = 14'b11111111111111;
	assign font[19][221] = 14'b11111111111111;
	assign font[20][221] = 14'b11111111111111;
	assign font[21][221] = 14'b11111111111111;
	assign font[22][221] = 14'b11111111111111;
	assign font[23][221] = 14'b11111111111111;
	assign font[24][221] = 14'b11111111111111;
	assign font[25][221] = 14'b11111111111111;
	assign font[26][221] = 14'b11111111111111;
	assign font[27][221] = 14'b11111111111111;
	assign font[28][221] = 14'b11111111111111;
	assign font[29][221] = 14'b11111111111111;
	assign font[30][221] = 14'b11111111111111;
	assign font[31][221] = 14'b11111111111111;

	assign font[0][222] = 14'b11111111111111;
	assign font[1][222] = 14'b11111111111111;
	assign font[2][222] = 14'b11111111111111;
	assign font[3][222] = 14'b11111111111111;
	assign font[4][222] = 14'b11111111111111;
	assign font[5][222] = 14'b11111111111111;
	assign font[6][222] = 14'b11111111111111;
	assign font[7][222] = 14'b11111111111111;
	assign font[8][222] = 14'b11111111111111;
	assign font[9][222] = 14'b11111111111111;
	assign font[10][222] = 14'b11111111111111;
	assign font[11][222] = 14'b11111111111111;
	assign font[12][222] = 14'b11111111111111;
	assign font[13][222] = 14'b11111111111111;
	assign font[14][222] = 14'b11111111111111;
	assign font[15][222] = 14'b11111111111111;
	assign font[16][222] = 14'b11111111111111;
	assign font[17][222] = 14'b11111111111111;
	assign font[18][222] = 14'b11111111111111;
	assign font[19][222] = 14'b11111111111111;
	assign font[20][222] = 14'b11111111111111;
	assign font[21][222] = 14'b11111111111111;
	assign font[22][222] = 14'b11111111111111;
	assign font[23][222] = 14'b11111111111111;
	assign font[24][222] = 14'b11111111111111;
	assign font[25][222] = 14'b11111111111111;
	assign font[26][222] = 14'b11111111111111;
	assign font[27][222] = 14'b11111111111111;
	assign font[28][222] = 14'b11111111111111;
	assign font[29][222] = 14'b11111111111111;
	assign font[30][222] = 14'b11111111111111;
	assign font[31][222] = 14'b11111111111111;

	assign font[0][223] = 14'b11111111111111;
	assign font[1][223] = 14'b11111111111111;
	assign font[2][223] = 14'b11111111111111;
	assign font[3][223] = 14'b11111111111111;
	assign font[4][223] = 14'b11111111111111;
	assign font[5][223] = 14'b11111111111111;
	assign font[6][223] = 14'b11111111111111;
	assign font[7][223] = 14'b11111111111111;
	assign font[8][223] = 14'b11111111111111;
	assign font[9][223] = 14'b11111111111111;
	assign font[10][223] = 14'b11111111111111;
	assign font[11][223] = 14'b11111111111111;
	assign font[12][223] = 14'b11111111111111;
	assign font[13][223] = 14'b11111111111111;
	assign font[14][223] = 14'b11111111111111;
	assign font[15][223] = 14'b11111111111111;
	assign font[16][223] = 14'b11111111111111;
	assign font[17][223] = 14'b11111111111111;
	assign font[18][223] = 14'b11111111111111;
	assign font[19][223] = 14'b11111111111111;
	assign font[20][223] = 14'b11111111111111;
	assign font[21][223] = 14'b11111111111111;
	assign font[22][223] = 14'b11111111111111;
	assign font[23][223] = 14'b11111111111111;
	assign font[24][223] = 14'b11111111111111;
	assign font[25][223] = 14'b11111111111111;
	assign font[26][223] = 14'b11111111111111;
	assign font[27][223] = 14'b11111111111111;
	assign font[28][223] = 14'b11111111111111;
	assign font[29][223] = 14'b11111111111111;
	assign font[30][223] = 14'b11111111111111;
	assign font[31][223] = 14'b11111111111111;

	assign font[0][224] = 14'b11111111111111;
	assign font[1][224] = 14'b11111111111111;
	assign font[2][224] = 14'b11111111111111;
	assign font[3][224] = 14'b11111111111111;
	assign font[4][224] = 14'b11111111111111;
	assign font[5][224] = 14'b11111111111111;
	assign font[6][224] = 14'b11111111111111;
	assign font[7][224] = 14'b11111111111111;
	assign font[8][224] = 14'b11111111111111;
	assign font[9][224] = 14'b11111111111111;
	assign font[10][224] = 14'b11111111111111;
	assign font[11][224] = 14'b11111111111111;
	assign font[12][224] = 14'b11111111111111;
	assign font[13][224] = 14'b11111111111111;
	assign font[14][224] = 14'b11111111111111;
	assign font[15][224] = 14'b11111111111111;
	assign font[16][224] = 14'b11111111111111;
	assign font[17][224] = 14'b11111111111111;
	assign font[18][224] = 14'b11111111111111;
	assign font[19][224] = 14'b11111111111111;
	assign font[20][224] = 14'b11111111111111;
	assign font[21][224] = 14'b11111111111111;
	assign font[22][224] = 14'b11111111111111;
	assign font[23][224] = 14'b11111111111111;
	assign font[24][224] = 14'b11111111111111;
	assign font[25][224] = 14'b11111111111111;
	assign font[26][224] = 14'b11111111111111;
	assign font[27][224] = 14'b11111111111111;
	assign font[28][224] = 14'b11111111111111;
	assign font[29][224] = 14'b11111111111111;
	assign font[30][224] = 14'b11111111111111;
	assign font[31][224] = 14'b11111111111111;

	assign font[0][225] = 14'b11111111111111;
	assign font[1][225] = 14'b11111111111111;
	assign font[2][225] = 14'b11111111111111;
	assign font[3][225] = 14'b11111111111111;
	assign font[4][225] = 14'b11111111111111;
	assign font[5][225] = 14'b11111111111111;
	assign font[6][225] = 14'b11111111111111;
	assign font[7][225] = 14'b11111111111111;
	assign font[8][225] = 14'b11111111111111;
	assign font[9][225] = 14'b11111111111111;
	assign font[10][225] = 14'b11111111111111;
	assign font[11][225] = 14'b11111111111111;
	assign font[12][225] = 14'b11111111111111;
	assign font[13][225] = 14'b11111111111111;
	assign font[14][225] = 14'b11111111111111;
	assign font[15][225] = 14'b11111111111111;
	assign font[16][225] = 14'b11111111111111;
	assign font[17][225] = 14'b11111111111111;
	assign font[18][225] = 14'b11111111111111;
	assign font[19][225] = 14'b11111111111111;
	assign font[20][225] = 14'b11111111111111;
	assign font[21][225] = 14'b11111111111111;
	assign font[22][225] = 14'b11111111111111;
	assign font[23][225] = 14'b11111111111111;
	assign font[24][225] = 14'b11111111111111;
	assign font[25][225] = 14'b11111111111111;
	assign font[26][225] = 14'b11111111111111;
	assign font[27][225] = 14'b11111111111111;
	assign font[28][225] = 14'b11111111111111;
	assign font[29][225] = 14'b11111111111111;
	assign font[30][225] = 14'b11111111111111;
	assign font[31][225] = 14'b11111111111111;

	assign font[0][226] = 14'b11111111111111;
	assign font[1][226] = 14'b11111111111111;
	assign font[2][226] = 14'b11111111111111;
	assign font[3][226] = 14'b11111111111111;
	assign font[4][226] = 14'b11111111111111;
	assign font[5][226] = 14'b11111111111111;
	assign font[6][226] = 14'b11111111111111;
	assign font[7][226] = 14'b11111111111111;
	assign font[8][226] = 14'b11111111111111;
	assign font[9][226] = 14'b11111111111111;
	assign font[10][226] = 14'b11111111111111;
	assign font[11][226] = 14'b11111111111111;
	assign font[12][226] = 14'b11111111111111;
	assign font[13][226] = 14'b11111111111111;
	assign font[14][226] = 14'b11111111111111;
	assign font[15][226] = 14'b11111111111111;
	assign font[16][226] = 14'b11111111111111;
	assign font[17][226] = 14'b11111111111111;
	assign font[18][226] = 14'b11111111111111;
	assign font[19][226] = 14'b11111111111111;
	assign font[20][226] = 14'b11111111111111;
	assign font[21][226] = 14'b11111111111111;
	assign font[22][226] = 14'b11111111111111;
	assign font[23][226] = 14'b11111111111111;
	assign font[24][226] = 14'b11111111111111;
	assign font[25][226] = 14'b11111111111111;
	assign font[26][226] = 14'b11111111111111;
	assign font[27][226] = 14'b11111111111111;
	assign font[28][226] = 14'b11111111111111;
	assign font[29][226] = 14'b11111111111111;
	assign font[30][226] = 14'b11111111111111;
	assign font[31][226] = 14'b11111111111111;

	assign font[0][227] = 14'b11111111111111;
	assign font[1][227] = 14'b11111111111111;
	assign font[2][227] = 14'b11111111111111;
	assign font[3][227] = 14'b11111111111111;
	assign font[4][227] = 14'b11111111111111;
	assign font[5][227] = 14'b11111111111111;
	assign font[6][227] = 14'b11111111111111;
	assign font[7][227] = 14'b11111111111111;
	assign font[8][227] = 14'b11111111111111;
	assign font[9][227] = 14'b11111111111111;
	assign font[10][227] = 14'b11111111111111;
	assign font[11][227] = 14'b11111111111111;
	assign font[12][227] = 14'b11111111111111;
	assign font[13][227] = 14'b11111111111111;
	assign font[14][227] = 14'b11111111111111;
	assign font[15][227] = 14'b11111111111111;
	assign font[16][227] = 14'b11111111111111;
	assign font[17][227] = 14'b11111111111111;
	assign font[18][227] = 14'b11111111111111;
	assign font[19][227] = 14'b11111111111111;
	assign font[20][227] = 14'b11111111111111;
	assign font[21][227] = 14'b11111111111111;
	assign font[22][227] = 14'b11111111111111;
	assign font[23][227] = 14'b11111111111111;
	assign font[24][227] = 14'b11111111111111;
	assign font[25][227] = 14'b11111111111111;
	assign font[26][227] = 14'b11111111111111;
	assign font[27][227] = 14'b11111111111111;
	assign font[28][227] = 14'b11111111111111;
	assign font[29][227] = 14'b11111111111111;
	assign font[30][227] = 14'b11111111111111;
	assign font[31][227] = 14'b11111111111111;

	assign font[0][228] = 14'b11111111111111;
	assign font[1][228] = 14'b11111111111111;
	assign font[2][228] = 14'b11111111111111;
	assign font[3][228] = 14'b11111111111111;
	assign font[4][228] = 14'b11111111111111;
	assign font[5][228] = 14'b11111111111111;
	assign font[6][228] = 14'b11111111111111;
	assign font[7][228] = 14'b11111111111111;
	assign font[8][228] = 14'b11111111111111;
	assign font[9][228] = 14'b11111111111111;
	assign font[10][228] = 14'b11111111111111;
	assign font[11][228] = 14'b11111111111111;
	assign font[12][228] = 14'b11111111111111;
	assign font[13][228] = 14'b11111111111111;
	assign font[14][228] = 14'b11111111111111;
	assign font[15][228] = 14'b11111111111111;
	assign font[16][228] = 14'b11111111111111;
	assign font[17][228] = 14'b11111111111111;
	assign font[18][228] = 14'b11111111111111;
	assign font[19][228] = 14'b11111111111111;
	assign font[20][228] = 14'b11111111111111;
	assign font[21][228] = 14'b11111111111111;
	assign font[22][228] = 14'b11111111111111;
	assign font[23][228] = 14'b11111111111111;
	assign font[24][228] = 14'b11111111111111;
	assign font[25][228] = 14'b11111111111111;
	assign font[26][228] = 14'b11111111111111;
	assign font[27][228] = 14'b11111111111111;
	assign font[28][228] = 14'b11111111111111;
	assign font[29][228] = 14'b11111111111111;
	assign font[30][228] = 14'b11111111111111;
	assign font[31][228] = 14'b11111111111111;

	assign font[0][229] = 14'b11111111111111;
	assign font[1][229] = 14'b11111111111111;
	assign font[2][229] = 14'b11111111111111;
	assign font[3][229] = 14'b11111111111111;
	assign font[4][229] = 14'b11111111111111;
	assign font[5][229] = 14'b11111111111111;
	assign font[6][229] = 14'b11111111111111;
	assign font[7][229] = 14'b11111111111111;
	assign font[8][229] = 14'b11111111111111;
	assign font[9][229] = 14'b11111111111111;
	assign font[10][229] = 14'b11111111111111;
	assign font[11][229] = 14'b11111111111111;
	assign font[12][229] = 14'b11111111111111;
	assign font[13][229] = 14'b11111111111111;
	assign font[14][229] = 14'b11111111111111;
	assign font[15][229] = 14'b11111111111111;
	assign font[16][229] = 14'b11111111111111;
	assign font[17][229] = 14'b11111111111111;
	assign font[18][229] = 14'b11111111111111;
	assign font[19][229] = 14'b11111111111111;
	assign font[20][229] = 14'b11111111111111;
	assign font[21][229] = 14'b11111111111111;
	assign font[22][229] = 14'b11111111111111;
	assign font[23][229] = 14'b11111111111111;
	assign font[24][229] = 14'b11111111111111;
	assign font[25][229] = 14'b11111111111111;
	assign font[26][229] = 14'b11111111111111;
	assign font[27][229] = 14'b11111111111111;
	assign font[28][229] = 14'b11111111111111;
	assign font[29][229] = 14'b11111111111111;
	assign font[30][229] = 14'b11111111111111;
	assign font[31][229] = 14'b11111111111111;

	assign font[0][230] = 14'b11111111111111;
	assign font[1][230] = 14'b11111111111111;
	assign font[2][230] = 14'b11111111111111;
	assign font[3][230] = 14'b11111111111111;
	assign font[4][230] = 14'b11111111111111;
	assign font[5][230] = 14'b11111111111111;
	assign font[6][230] = 14'b11111111111111;
	assign font[7][230] = 14'b11111111111111;
	assign font[8][230] = 14'b11111111111111;
	assign font[9][230] = 14'b11111111111111;
	assign font[10][230] = 14'b11111111111111;
	assign font[11][230] = 14'b11111111111111;
	assign font[12][230] = 14'b11111111111111;
	assign font[13][230] = 14'b11111111111111;
	assign font[14][230] = 14'b11111111111111;
	assign font[15][230] = 14'b11111111111111;
	assign font[16][230] = 14'b11111111111111;
	assign font[17][230] = 14'b11111111111111;
	assign font[18][230] = 14'b11111111111111;
	assign font[19][230] = 14'b11111111111111;
	assign font[20][230] = 14'b11111111111111;
	assign font[21][230] = 14'b11111111111111;
	assign font[22][230] = 14'b11111111111111;
	assign font[23][230] = 14'b11111111111111;
	assign font[24][230] = 14'b11111111111111;
	assign font[25][230] = 14'b11111111111111;
	assign font[26][230] = 14'b11111111111111;
	assign font[27][230] = 14'b11111111111111;
	assign font[28][230] = 14'b11111111111111;
	assign font[29][230] = 14'b11111111111111;
	assign font[30][230] = 14'b11111111111111;
	assign font[31][230] = 14'b11111111111111;

	assign font[0][231] = 14'b11111111111111;
	assign font[1][231] = 14'b11111111111111;
	assign font[2][231] = 14'b11111111111111;
	assign font[3][231] = 14'b11111111111111;
	assign font[4][231] = 14'b11111111111111;
	assign font[5][231] = 14'b11111111111111;
	assign font[6][231] = 14'b11111111111111;
	assign font[7][231] = 14'b11111111111111;
	assign font[8][231] = 14'b11111111111111;
	assign font[9][231] = 14'b11111111111111;
	assign font[10][231] = 14'b11111111111111;
	assign font[11][231] = 14'b11111111111111;
	assign font[12][231] = 14'b11111111111111;
	assign font[13][231] = 14'b11111111111111;
	assign font[14][231] = 14'b11111111111111;
	assign font[15][231] = 14'b11111111111111;
	assign font[16][231] = 14'b11111111111111;
	assign font[17][231] = 14'b11111111111111;
	assign font[18][231] = 14'b11111111111111;
	assign font[19][231] = 14'b11111111111111;
	assign font[20][231] = 14'b11111111111111;
	assign font[21][231] = 14'b11111111111111;
	assign font[22][231] = 14'b11111111111111;
	assign font[23][231] = 14'b11111111111111;
	assign font[24][231] = 14'b11111111111111;
	assign font[25][231] = 14'b11111111111111;
	assign font[26][231] = 14'b11111111111111;
	assign font[27][231] = 14'b11111111111111;
	assign font[28][231] = 14'b11111111111111;
	assign font[29][231] = 14'b11111111111111;
	assign font[30][231] = 14'b11111111111111;
	assign font[31][231] = 14'b11111111111111;

	assign font[0][232] = 14'b11111111111111;
	assign font[1][232] = 14'b11111111111111;
	assign font[2][232] = 14'b11111111111111;
	assign font[3][232] = 14'b11111111111111;
	assign font[4][232] = 14'b11111111111111;
	assign font[5][232] = 14'b11111111111111;
	assign font[6][232] = 14'b11111111111111;
	assign font[7][232] = 14'b11111111111111;
	assign font[8][232] = 14'b11111111111111;
	assign font[9][232] = 14'b11111111111111;
	assign font[10][232] = 14'b11111111111111;
	assign font[11][232] = 14'b11111111111111;
	assign font[12][232] = 14'b11111111111111;
	assign font[13][232] = 14'b11111111111111;
	assign font[14][232] = 14'b11111111111111;
	assign font[15][232] = 14'b11111111111111;
	assign font[16][232] = 14'b11111111111111;
	assign font[17][232] = 14'b11111111111111;
	assign font[18][232] = 14'b11111111111111;
	assign font[19][232] = 14'b11111111111111;
	assign font[20][232] = 14'b11111111111111;
	assign font[21][232] = 14'b11111111111111;
	assign font[22][232] = 14'b11111111111111;
	assign font[23][232] = 14'b11111111111111;
	assign font[24][232] = 14'b11111111111111;
	assign font[25][232] = 14'b11111111111111;
	assign font[26][232] = 14'b11111111111111;
	assign font[27][232] = 14'b11111111111111;
	assign font[28][232] = 14'b11111111111111;
	assign font[29][232] = 14'b11111111111111;
	assign font[30][232] = 14'b11111111111111;
	assign font[31][232] = 14'b11111111111111;

	assign font[0][233] = 14'b11111111111111;
	assign font[1][233] = 14'b11111111111111;
	assign font[2][233] = 14'b11111111111111;
	assign font[3][233] = 14'b11111111111111;
	assign font[4][233] = 14'b11111111111111;
	assign font[5][233] = 14'b11111111111111;
	assign font[6][233] = 14'b11111111111111;
	assign font[7][233] = 14'b11111111111111;
	assign font[8][233] = 14'b11111111111111;
	assign font[9][233] = 14'b11111111111111;
	assign font[10][233] = 14'b11111111111111;
	assign font[11][233] = 14'b11111111111111;
	assign font[12][233] = 14'b11111111111111;
	assign font[13][233] = 14'b11111111111111;
	assign font[14][233] = 14'b11111111111111;
	assign font[15][233] = 14'b11111111111111;
	assign font[16][233] = 14'b11111111111111;
	assign font[17][233] = 14'b11111111111111;
	assign font[18][233] = 14'b11111111111111;
	assign font[19][233] = 14'b11111111111111;
	assign font[20][233] = 14'b11111111111111;
	assign font[21][233] = 14'b11111111111111;
	assign font[22][233] = 14'b11111111111111;
	assign font[23][233] = 14'b11111111111111;
	assign font[24][233] = 14'b11111111111111;
	assign font[25][233] = 14'b11111111111111;
	assign font[26][233] = 14'b11111111111111;
	assign font[27][233] = 14'b11111111111111;
	assign font[28][233] = 14'b11111111111111;
	assign font[29][233] = 14'b11111111111111;
	assign font[30][233] = 14'b11111111111111;
	assign font[31][233] = 14'b11111111111111;

	assign font[0][234] = 14'b11111111111111;
	assign font[1][234] = 14'b11111111111111;
	assign font[2][234] = 14'b11111111111111;
	assign font[3][234] = 14'b11111111111111;
	assign font[4][234] = 14'b11111111111111;
	assign font[5][234] = 14'b11111111111111;
	assign font[6][234] = 14'b11111111111111;
	assign font[7][234] = 14'b11111111111111;
	assign font[8][234] = 14'b11111111111111;
	assign font[9][234] = 14'b11111111111111;
	assign font[10][234] = 14'b11111111111111;
	assign font[11][234] = 14'b11111111111111;
	assign font[12][234] = 14'b11111111111111;
	assign font[13][234] = 14'b11111111111111;
	assign font[14][234] = 14'b11111111111111;
	assign font[15][234] = 14'b11111111111111;
	assign font[16][234] = 14'b11111111111111;
	assign font[17][234] = 14'b11111111111111;
	assign font[18][234] = 14'b11111111111111;
	assign font[19][234] = 14'b11111111111111;
	assign font[20][234] = 14'b11111111111111;
	assign font[21][234] = 14'b11111111111111;
	assign font[22][234] = 14'b11111111111111;
	assign font[23][234] = 14'b11111111111111;
	assign font[24][234] = 14'b11111111111111;
	assign font[25][234] = 14'b11111111111111;
	assign font[26][234] = 14'b11111111111111;
	assign font[27][234] = 14'b11111111111111;
	assign font[28][234] = 14'b11111111111111;
	assign font[29][234] = 14'b11111111111111;
	assign font[30][234] = 14'b11111111111111;
	assign font[31][234] = 14'b11111111111111;

	assign font[0][235] = 14'b11111111111111;
	assign font[1][235] = 14'b11111111111111;
	assign font[2][235] = 14'b11111111111111;
	assign font[3][235] = 14'b11111111111111;
	assign font[4][235] = 14'b11111111111111;
	assign font[5][235] = 14'b11111111111111;
	assign font[6][235] = 14'b11111111111111;
	assign font[7][235] = 14'b11111111111111;
	assign font[8][235] = 14'b11111111111111;
	assign font[9][235] = 14'b11111111111111;
	assign font[10][235] = 14'b11111111111111;
	assign font[11][235] = 14'b11111111111111;
	assign font[12][235] = 14'b11111111111111;
	assign font[13][235] = 14'b11111111111111;
	assign font[14][235] = 14'b11111111111111;
	assign font[15][235] = 14'b11111111111111;
	assign font[16][235] = 14'b11111111111111;
	assign font[17][235] = 14'b11111111111111;
	assign font[18][235] = 14'b11111111111111;
	assign font[19][235] = 14'b11111111111111;
	assign font[20][235] = 14'b11111111111111;
	assign font[21][235] = 14'b11111111111111;
	assign font[22][235] = 14'b11111111111111;
	assign font[23][235] = 14'b11111111111111;
	assign font[24][235] = 14'b11111111111111;
	assign font[25][235] = 14'b11111111111111;
	assign font[26][235] = 14'b11111111111111;
	assign font[27][235] = 14'b11111111111111;
	assign font[28][235] = 14'b11111111111111;
	assign font[29][235] = 14'b11111111111111;
	assign font[30][235] = 14'b11111111111111;
	assign font[31][235] = 14'b11111111111111;

	assign font[0][236] = 14'b11111111111111;
	assign font[1][236] = 14'b11111111111111;
	assign font[2][236] = 14'b11111111111111;
	assign font[3][236] = 14'b11111111111111;
	assign font[4][236] = 14'b11111111111111;
	assign font[5][236] = 14'b11111111111111;
	assign font[6][236] = 14'b11111111111111;
	assign font[7][236] = 14'b11111111111111;
	assign font[8][236] = 14'b11111111111111;
	assign font[9][236] = 14'b11111111111111;
	assign font[10][236] = 14'b11111111111111;
	assign font[11][236] = 14'b11111111111111;
	assign font[12][236] = 14'b11111111111111;
	assign font[13][236] = 14'b11111111111111;
	assign font[14][236] = 14'b11111111111111;
	assign font[15][236] = 14'b11111111111111;
	assign font[16][236] = 14'b11111111111111;
	assign font[17][236] = 14'b11111111111111;
	assign font[18][236] = 14'b11111111111111;
	assign font[19][236] = 14'b11111111111111;
	assign font[20][236] = 14'b11111111111111;
	assign font[21][236] = 14'b11111111111111;
	assign font[22][236] = 14'b11111111111111;
	assign font[23][236] = 14'b11111111111111;
	assign font[24][236] = 14'b11111111111111;
	assign font[25][236] = 14'b11111111111111;
	assign font[26][236] = 14'b11111111111111;
	assign font[27][236] = 14'b11111111111111;
	assign font[28][236] = 14'b11111111111111;
	assign font[29][236] = 14'b11111111111111;
	assign font[30][236] = 14'b11111111111111;
	assign font[31][236] = 14'b11111111111111;

	assign font[0][237] = 14'b11111111111111;
	assign font[1][237] = 14'b11111111111111;
	assign font[2][237] = 14'b11111111111111;
	assign font[3][237] = 14'b11111111111111;
	assign font[4][237] = 14'b11111111111111;
	assign font[5][237] = 14'b11111111111111;
	assign font[6][237] = 14'b11111111111111;
	assign font[7][237] = 14'b11111111111111;
	assign font[8][237] = 14'b11111111111111;
	assign font[9][237] = 14'b11111111111111;
	assign font[10][237] = 14'b11111111111111;
	assign font[11][237] = 14'b11111111111111;
	assign font[12][237] = 14'b11111111111111;
	assign font[13][237] = 14'b11111111111111;
	assign font[14][237] = 14'b11111111111111;
	assign font[15][237] = 14'b11111111111111;
	assign font[16][237] = 14'b11111111111111;
	assign font[17][237] = 14'b11111111111111;
	assign font[18][237] = 14'b11111111111111;
	assign font[19][237] = 14'b11111111111111;
	assign font[20][237] = 14'b11111111111111;
	assign font[21][237] = 14'b11111111111111;
	assign font[22][237] = 14'b11111111111111;
	assign font[23][237] = 14'b11111111111111;
	assign font[24][237] = 14'b11111111111111;
	assign font[25][237] = 14'b11111111111111;
	assign font[26][237] = 14'b11111111111111;
	assign font[27][237] = 14'b11111111111111;
	assign font[28][237] = 14'b11111111111111;
	assign font[29][237] = 14'b11111111111111;
	assign font[30][237] = 14'b11111111111111;
	assign font[31][237] = 14'b11111111111111;

	assign font[0][238] = 14'b11111111111111;
	assign font[1][238] = 14'b11111111111111;
	assign font[2][238] = 14'b11111111111111;
	assign font[3][238] = 14'b11111111111111;
	assign font[4][238] = 14'b11111111111111;
	assign font[5][238] = 14'b11111111111111;
	assign font[6][238] = 14'b11111111111111;
	assign font[7][238] = 14'b11111111111111;
	assign font[8][238] = 14'b11111111111111;
	assign font[9][238] = 14'b11111111111111;
	assign font[10][238] = 14'b11111111111111;
	assign font[11][238] = 14'b11111111111111;
	assign font[12][238] = 14'b11111111111111;
	assign font[13][238] = 14'b11111111111111;
	assign font[14][238] = 14'b11111111111111;
	assign font[15][238] = 14'b11111111111111;
	assign font[16][238] = 14'b11111111111111;
	assign font[17][238] = 14'b11111111111111;
	assign font[18][238] = 14'b11111111111111;
	assign font[19][238] = 14'b11111111111111;
	assign font[20][238] = 14'b11111111111111;
	assign font[21][238] = 14'b11111111111111;
	assign font[22][238] = 14'b11111111111111;
	assign font[23][238] = 14'b11111111111111;
	assign font[24][238] = 14'b11111111111111;
	assign font[25][238] = 14'b11111111111111;
	assign font[26][238] = 14'b11111111111111;
	assign font[27][238] = 14'b11111111111111;
	assign font[28][238] = 14'b11111111111111;
	assign font[29][238] = 14'b11111111111111;
	assign font[30][238] = 14'b11111111111111;
	assign font[31][238] = 14'b11111111111111;

	assign font[0][239] = 14'b11111111111111;
	assign font[1][239] = 14'b11111111111111;
	assign font[2][239] = 14'b11111111111111;
	assign font[3][239] = 14'b11111111111111;
	assign font[4][239] = 14'b11111111111111;
	assign font[5][239] = 14'b11111111111111;
	assign font[6][239] = 14'b11111111111111;
	assign font[7][239] = 14'b11111111111111;
	assign font[8][239] = 14'b11111111111111;
	assign font[9][239] = 14'b11111111111111;
	assign font[10][239] = 14'b11111111111111;
	assign font[11][239] = 14'b11111111111111;
	assign font[12][239] = 14'b11111111111111;
	assign font[13][239] = 14'b11111111111111;
	assign font[14][239] = 14'b11111111111111;
	assign font[15][239] = 14'b11111111111111;
	assign font[16][239] = 14'b11111111111111;
	assign font[17][239] = 14'b11111111111111;
	assign font[18][239] = 14'b11111111111111;
	assign font[19][239] = 14'b11111111111111;
	assign font[20][239] = 14'b11111111111111;
	assign font[21][239] = 14'b11111111111111;
	assign font[22][239] = 14'b11111111111111;
	assign font[23][239] = 14'b11111111111111;
	assign font[24][239] = 14'b11111111111111;
	assign font[25][239] = 14'b11111111111111;
	assign font[26][239] = 14'b11111111111111;
	assign font[27][239] = 14'b11111111111111;
	assign font[28][239] = 14'b11111111111111;
	assign font[29][239] = 14'b11111111111111;
	assign font[30][239] = 14'b11111111111111;
	assign font[31][239] = 14'b11111111111111;

	assign font[0][240] = 14'b11111111111111;
	assign font[1][240] = 14'b11111111111111;
	assign font[2][240] = 14'b11111111111111;
	assign font[3][240] = 14'b11111111111111;
	assign font[4][240] = 14'b11111111111111;
	assign font[5][240] = 14'b11111111111111;
	assign font[6][240] = 14'b11111111111111;
	assign font[7][240] = 14'b11111111111111;
	assign font[8][240] = 14'b11111111111111;
	assign font[9][240] = 14'b11111111111111;
	assign font[10][240] = 14'b11111111111111;
	assign font[11][240] = 14'b11111111111111;
	assign font[12][240] = 14'b11111111111111;
	assign font[13][240] = 14'b11111111111111;
	assign font[14][240] = 14'b11111111111111;
	assign font[15][240] = 14'b11111111111111;
	assign font[16][240] = 14'b11111111111111;
	assign font[17][240] = 14'b11111111111111;
	assign font[18][240] = 14'b11111111111111;
	assign font[19][240] = 14'b11111111111111;
	assign font[20][240] = 14'b11111111111111;
	assign font[21][240] = 14'b11111111111111;
	assign font[22][240] = 14'b11111111111111;
	assign font[23][240] = 14'b11111111111111;
	assign font[24][240] = 14'b11111111111111;
	assign font[25][240] = 14'b11111111111111;
	assign font[26][240] = 14'b11111111111111;
	assign font[27][240] = 14'b11111111111111;
	assign font[28][240] = 14'b11111111111111;
	assign font[29][240] = 14'b11111111111111;
	assign font[30][240] = 14'b11111111111111;
	assign font[31][240] = 14'b11111111111111;

	assign font[0][241] = 14'b11111111111111;
	assign font[1][241] = 14'b11111111111111;
	assign font[2][241] = 14'b11111111111111;
	assign font[3][241] = 14'b11111111111111;
	assign font[4][241] = 14'b11111111111111;
	assign font[5][241] = 14'b11111111111111;
	assign font[6][241] = 14'b11111111111111;
	assign font[7][241] = 14'b11111111111111;
	assign font[8][241] = 14'b11111111111111;
	assign font[9][241] = 14'b11111111111111;
	assign font[10][241] = 14'b11111111111111;
	assign font[11][241] = 14'b11111111111111;
	assign font[12][241] = 14'b11111111111111;
	assign font[13][241] = 14'b11111111111111;
	assign font[14][241] = 14'b11111111111111;
	assign font[15][241] = 14'b11111111111111;
	assign font[16][241] = 14'b11111111111111;
	assign font[17][241] = 14'b11111111111111;
	assign font[18][241] = 14'b11111111111111;
	assign font[19][241] = 14'b11111111111111;
	assign font[20][241] = 14'b11111111111111;
	assign font[21][241] = 14'b11111111111111;
	assign font[22][241] = 14'b11111111111111;
	assign font[23][241] = 14'b11111111111111;
	assign font[24][241] = 14'b11111111111111;
	assign font[25][241] = 14'b11111111111111;
	assign font[26][241] = 14'b11111111111111;
	assign font[27][241] = 14'b11111111111111;
	assign font[28][241] = 14'b11111111111111;
	assign font[29][241] = 14'b11111111111111;
	assign font[30][241] = 14'b11111111111111;
	assign font[31][241] = 14'b11111111111111;

	assign font[0][242] = 14'b11111111111111;
	assign font[1][242] = 14'b11111111111111;
	assign font[2][242] = 14'b11111111111111;
	assign font[3][242] = 14'b11111111111111;
	assign font[4][242] = 14'b11111111111111;
	assign font[5][242] = 14'b11111111111111;
	assign font[6][242] = 14'b11111111111111;
	assign font[7][242] = 14'b11111111111111;
	assign font[8][242] = 14'b11111111111111;
	assign font[9][242] = 14'b11111111111111;
	assign font[10][242] = 14'b11111111111111;
	assign font[11][242] = 14'b11111111111111;
	assign font[12][242] = 14'b11111111111111;
	assign font[13][242] = 14'b11111111111111;
	assign font[14][242] = 14'b11111111111111;
	assign font[15][242] = 14'b11111111111111;
	assign font[16][242] = 14'b11111111111111;
	assign font[17][242] = 14'b11111111111111;
	assign font[18][242] = 14'b11111111111111;
	assign font[19][242] = 14'b11111111111111;
	assign font[20][242] = 14'b11111111111111;
	assign font[21][242] = 14'b11111111111111;
	assign font[22][242] = 14'b11111111111111;
	assign font[23][242] = 14'b11111111111111;
	assign font[24][242] = 14'b11111111111111;
	assign font[25][242] = 14'b11111111111111;
	assign font[26][242] = 14'b11111111111111;
	assign font[27][242] = 14'b11111111111111;
	assign font[28][242] = 14'b11111111111111;
	assign font[29][242] = 14'b11111111111111;
	assign font[30][242] = 14'b11111111111111;
	assign font[31][242] = 14'b11111111111111;

	assign font[0][243] = 14'b11111111111111;
	assign font[1][243] = 14'b11111111111111;
	assign font[2][243] = 14'b11111111111111;
	assign font[3][243] = 14'b11111111111111;
	assign font[4][243] = 14'b11111111111111;
	assign font[5][243] = 14'b11111111111111;
	assign font[6][243] = 14'b11111111111111;
	assign font[7][243] = 14'b11111111111111;
	assign font[8][243] = 14'b11111111111111;
	assign font[9][243] = 14'b11111111111111;
	assign font[10][243] = 14'b11111111111111;
	assign font[11][243] = 14'b11111111111111;
	assign font[12][243] = 14'b11111111111111;
	assign font[13][243] = 14'b11111111111111;
	assign font[14][243] = 14'b11111111111111;
	assign font[15][243] = 14'b11111111111111;
	assign font[16][243] = 14'b11111111111111;
	assign font[17][243] = 14'b11111111111111;
	assign font[18][243] = 14'b11111111111111;
	assign font[19][243] = 14'b11111111111111;
	assign font[20][243] = 14'b11111111111111;
	assign font[21][243] = 14'b11111111111111;
	assign font[22][243] = 14'b11111111111111;
	assign font[23][243] = 14'b11111111111111;
	assign font[24][243] = 14'b11111111111111;
	assign font[25][243] = 14'b11111111111111;
	assign font[26][243] = 14'b11111111111111;
	assign font[27][243] = 14'b11111111111111;
	assign font[28][243] = 14'b11111111111111;
	assign font[29][243] = 14'b11111111111111;
	assign font[30][243] = 14'b11111111111111;
	assign font[31][243] = 14'b11111111111111;

	assign font[0][244] = 14'b11111111111111;
	assign font[1][244] = 14'b11111111111111;
	assign font[2][244] = 14'b11111111111111;
	assign font[3][244] = 14'b11111111111111;
	assign font[4][244] = 14'b11111111111111;
	assign font[5][244] = 14'b11111111111111;
	assign font[6][244] = 14'b11111111111111;
	assign font[7][244] = 14'b11111111111111;
	assign font[8][244] = 14'b11111111111111;
	assign font[9][244] = 14'b11111111111111;
	assign font[10][244] = 14'b11111111111111;
	assign font[11][244] = 14'b11111111111111;
	assign font[12][244] = 14'b11111111111111;
	assign font[13][244] = 14'b11111111111111;
	assign font[14][244] = 14'b11111111111111;
	assign font[15][244] = 14'b11111111111111;
	assign font[16][244] = 14'b11111111111111;
	assign font[17][244] = 14'b11111111111111;
	assign font[18][244] = 14'b11111111111111;
	assign font[19][244] = 14'b11111111111111;
	assign font[20][244] = 14'b11111111111111;
	assign font[21][244] = 14'b11111111111111;
	assign font[22][244] = 14'b11111111111111;
	assign font[23][244] = 14'b11111111111111;
	assign font[24][244] = 14'b11111111111111;
	assign font[25][244] = 14'b11111111111111;
	assign font[26][244] = 14'b11111111111111;
	assign font[27][244] = 14'b11111111111111;
	assign font[28][244] = 14'b11111111111111;
	assign font[29][244] = 14'b11111111111111;
	assign font[30][244] = 14'b11111111111111;
	assign font[31][244] = 14'b11111111111111;

	assign font[0][245] = 14'b11111111111111;
	assign font[1][245] = 14'b11111111111111;
	assign font[2][245] = 14'b11111111111111;
	assign font[3][245] = 14'b11111111111111;
	assign font[4][245] = 14'b11111111111111;
	assign font[5][245] = 14'b11111111111111;
	assign font[6][245] = 14'b11111111111111;
	assign font[7][245] = 14'b11111111111111;
	assign font[8][245] = 14'b11111111111111;
	assign font[9][245] = 14'b11111111111111;
	assign font[10][245] = 14'b11111111111111;
	assign font[11][245] = 14'b11111111111111;
	assign font[12][245] = 14'b11111111111111;
	assign font[13][245] = 14'b11111111111111;
	assign font[14][245] = 14'b11111111111111;
	assign font[15][245] = 14'b11111111111111;
	assign font[16][245] = 14'b11111111111111;
	assign font[17][245] = 14'b11111111111111;
	assign font[18][245] = 14'b11111111111111;
	assign font[19][245] = 14'b11111111111111;
	assign font[20][245] = 14'b11111111111111;
	assign font[21][245] = 14'b11111111111111;
	assign font[22][245] = 14'b11111111111111;
	assign font[23][245] = 14'b11111111111111;
	assign font[24][245] = 14'b11111111111111;
	assign font[25][245] = 14'b11111111111111;
	assign font[26][245] = 14'b11111111111111;
	assign font[27][245] = 14'b11111111111111;
	assign font[28][245] = 14'b11111111111111;
	assign font[29][245] = 14'b11111111111111;
	assign font[30][245] = 14'b11111111111111;
	assign font[31][245] = 14'b11111111111111;

	assign font[0][246] = 14'b11111111111111;
	assign font[1][246] = 14'b11111111111111;
	assign font[2][246] = 14'b11111111111111;
	assign font[3][246] = 14'b11111111111111;
	assign font[4][246] = 14'b11111111111111;
	assign font[5][246] = 14'b11111111111111;
	assign font[6][246] = 14'b11111111111111;
	assign font[7][246] = 14'b11111111111111;
	assign font[8][246] = 14'b11111111111111;
	assign font[9][246] = 14'b11111111111111;
	assign font[10][246] = 14'b11111111111111;
	assign font[11][246] = 14'b11111111111111;
	assign font[12][246] = 14'b11111111111111;
	assign font[13][246] = 14'b11111111111111;
	assign font[14][246] = 14'b11111111111111;
	assign font[15][246] = 14'b11111111111111;
	assign font[16][246] = 14'b11111111111111;
	assign font[17][246] = 14'b11111111111111;
	assign font[18][246] = 14'b11111111111111;
	assign font[19][246] = 14'b11111111111111;
	assign font[20][246] = 14'b11111111111111;
	assign font[21][246] = 14'b11111111111111;
	assign font[22][246] = 14'b11111111111111;
	assign font[23][246] = 14'b11111111111111;
	assign font[24][246] = 14'b11111111111111;
	assign font[25][246] = 14'b11111111111111;
	assign font[26][246] = 14'b11111111111111;
	assign font[27][246] = 14'b11111111111111;
	assign font[28][246] = 14'b11111111111111;
	assign font[29][246] = 14'b11111111111111;
	assign font[30][246] = 14'b11111111111111;
	assign font[31][246] = 14'b11111111111111;

	assign font[0][247] = 14'b11111111111111;
	assign font[1][247] = 14'b11111111111111;
	assign font[2][247] = 14'b11111111111111;
	assign font[3][247] = 14'b11111111111111;
	assign font[4][247] = 14'b11111111111111;
	assign font[5][247] = 14'b11111111111111;
	assign font[6][247] = 14'b11111111111111;
	assign font[7][247] = 14'b11111111111111;
	assign font[8][247] = 14'b11111111111111;
	assign font[9][247] = 14'b11111111111111;
	assign font[10][247] = 14'b11111111111111;
	assign font[11][247] = 14'b11111111111111;
	assign font[12][247] = 14'b11111111111111;
	assign font[13][247] = 14'b11111111111111;
	assign font[14][247] = 14'b11111111111111;
	assign font[15][247] = 14'b11111111111111;
	assign font[16][247] = 14'b11111111111111;
	assign font[17][247] = 14'b11111111111111;
	assign font[18][247] = 14'b11111111111111;
	assign font[19][247] = 14'b11111111111111;
	assign font[20][247] = 14'b11111111111111;
	assign font[21][247] = 14'b11111111111111;
	assign font[22][247] = 14'b11111111111111;
	assign font[23][247] = 14'b11111111111111;
	assign font[24][247] = 14'b11111111111111;
	assign font[25][247] = 14'b11111111111111;
	assign font[26][247] = 14'b11111111111111;
	assign font[27][247] = 14'b11111111111111;
	assign font[28][247] = 14'b11111111111111;
	assign font[29][247] = 14'b11111111111111;
	assign font[30][247] = 14'b11111111111111;
	assign font[31][247] = 14'b11111111111111;

	assign font[0][248] = 14'b11111111111111;
	assign font[1][248] = 14'b11111111111111;
	assign font[2][248] = 14'b11111111111111;
	assign font[3][248] = 14'b11111111111111;
	assign font[4][248] = 14'b11111111111111;
	assign font[5][248] = 14'b11111111111111;
	assign font[6][248] = 14'b11111111111111;
	assign font[7][248] = 14'b11111111111111;
	assign font[8][248] = 14'b11111111111111;
	assign font[9][248] = 14'b11111111111111;
	assign font[10][248] = 14'b11111111111111;
	assign font[11][248] = 14'b11111111111111;
	assign font[12][248] = 14'b11111111111111;
	assign font[13][248] = 14'b11111111111111;
	assign font[14][248] = 14'b11111111111111;
	assign font[15][248] = 14'b11111111111111;
	assign font[16][248] = 14'b11111111111111;
	assign font[17][248] = 14'b11111111111111;
	assign font[18][248] = 14'b11111111111111;
	assign font[19][248] = 14'b11111111111111;
	assign font[20][248] = 14'b11111111111111;
	assign font[21][248] = 14'b11111111111111;
	assign font[22][248] = 14'b11111111111111;
	assign font[23][248] = 14'b11111111111111;
	assign font[24][248] = 14'b11111111111111;
	assign font[25][248] = 14'b11111111111111;
	assign font[26][248] = 14'b11111111111111;
	assign font[27][248] = 14'b11111111111111;
	assign font[28][248] = 14'b11111111111111;
	assign font[29][248] = 14'b11111111111111;
	assign font[30][248] = 14'b11111111111111;
	assign font[31][248] = 14'b11111111111111;

	assign font[0][249] = 14'b11111111111111;
	assign font[1][249] = 14'b11111111111111;
	assign font[2][249] = 14'b11111111111111;
	assign font[3][249] = 14'b11111111111111;
	assign font[4][249] = 14'b11111111111111;
	assign font[5][249] = 14'b11111111111111;
	assign font[6][249] = 14'b11111111111111;
	assign font[7][249] = 14'b11111111111111;
	assign font[8][249] = 14'b11111111111111;
	assign font[9][249] = 14'b11111111111111;
	assign font[10][249] = 14'b11111111111111;
	assign font[11][249] = 14'b11111111111111;
	assign font[12][249] = 14'b11111111111111;
	assign font[13][249] = 14'b11111111111111;
	assign font[14][249] = 14'b11111111111111;
	assign font[15][249] = 14'b11111111111111;
	assign font[16][249] = 14'b11111111111111;
	assign font[17][249] = 14'b11111111111111;
	assign font[18][249] = 14'b11111111111111;
	assign font[19][249] = 14'b11111111111111;
	assign font[20][249] = 14'b11111111111111;
	assign font[21][249] = 14'b11111111111111;
	assign font[22][249] = 14'b11111111111111;
	assign font[23][249] = 14'b11111111111111;
	assign font[24][249] = 14'b11111111111111;
	assign font[25][249] = 14'b11111111111111;
	assign font[26][249] = 14'b11111111111111;
	assign font[27][249] = 14'b11111111111111;
	assign font[28][249] = 14'b11111111111111;
	assign font[29][249] = 14'b11111111111111;
	assign font[30][249] = 14'b11111111111111;
	assign font[31][249] = 14'b11111111111111;

	assign font[0][250] = 14'b11111111111111;
	assign font[1][250] = 14'b11111111111111;
	assign font[2][250] = 14'b11111111111111;
	assign font[3][250] = 14'b11111111111111;
	assign font[4][250] = 14'b11111111111111;
	assign font[5][250] = 14'b11111111111111;
	assign font[6][250] = 14'b11111111111111;
	assign font[7][250] = 14'b11111111111111;
	assign font[8][250] = 14'b11111111111111;
	assign font[9][250] = 14'b11111111111111;
	assign font[10][250] = 14'b11111111111111;
	assign font[11][250] = 14'b11111111111111;
	assign font[12][250] = 14'b11111111111111;
	assign font[13][250] = 14'b11111111111111;
	assign font[14][250] = 14'b11111111111111;
	assign font[15][250] = 14'b11111111111111;
	assign font[16][250] = 14'b11111111111111;
	assign font[17][250] = 14'b11111111111111;
	assign font[18][250] = 14'b11111111111111;
	assign font[19][250] = 14'b11111111111111;
	assign font[20][250] = 14'b11111111111111;
	assign font[21][250] = 14'b11111111111111;
	assign font[22][250] = 14'b11111111111111;
	assign font[23][250] = 14'b11111111111111;
	assign font[24][250] = 14'b11111111111111;
	assign font[25][250] = 14'b11111111111111;
	assign font[26][250] = 14'b11111111111111;
	assign font[27][250] = 14'b11111111111111;
	assign font[28][250] = 14'b11111111111111;
	assign font[29][250] = 14'b11111111111111;
	assign font[30][250] = 14'b11111111111111;
	assign font[31][250] = 14'b11111111111111;

	assign font[0][251] = 14'b11111111111111;
	assign font[1][251] = 14'b11111111111111;
	assign font[2][251] = 14'b11111111111111;
	assign font[3][251] = 14'b11111111111111;
	assign font[4][251] = 14'b11111111111111;
	assign font[5][251] = 14'b11111111111111;
	assign font[6][251] = 14'b11111111111111;
	assign font[7][251] = 14'b11111111111111;
	assign font[8][251] = 14'b11111111111111;
	assign font[9][251] = 14'b11111111111111;
	assign font[10][251] = 14'b11111111111111;
	assign font[11][251] = 14'b11111111111111;
	assign font[12][251] = 14'b11111111111111;
	assign font[13][251] = 14'b11111111111111;
	assign font[14][251] = 14'b11111111111111;
	assign font[15][251] = 14'b11111111111111;
	assign font[16][251] = 14'b11111111111111;
	assign font[17][251] = 14'b11111111111111;
	assign font[18][251] = 14'b11111111111111;
	assign font[19][251] = 14'b11111111111111;
	assign font[20][251] = 14'b11111111111111;
	assign font[21][251] = 14'b11111111111111;
	assign font[22][251] = 14'b11111111111111;
	assign font[23][251] = 14'b11111111111111;
	assign font[24][251] = 14'b11111111111111;
	assign font[25][251] = 14'b11111111111111;
	assign font[26][251] = 14'b11111111111111;
	assign font[27][251] = 14'b11111111111111;
	assign font[28][251] = 14'b11111111111111;
	assign font[29][251] = 14'b11111111111111;
	assign font[30][251] = 14'b11111111111111;
	assign font[31][251] = 14'b11111111111111;

	assign font[0][252] = 14'b11111111111111;
	assign font[1][252] = 14'b11111111111111;
	assign font[2][252] = 14'b11111111111111;
	assign font[3][252] = 14'b11111111111111;
	assign font[4][252] = 14'b11111111111111;
	assign font[5][252] = 14'b11111111111111;
	assign font[6][252] = 14'b11111111111111;
	assign font[7][252] = 14'b11111111111111;
	assign font[8][252] = 14'b11111111111111;
	assign font[9][252] = 14'b11111111111111;
	assign font[10][252] = 14'b11111111111111;
	assign font[11][252] = 14'b11111111111111;
	assign font[12][252] = 14'b11111111111111;
	assign font[13][252] = 14'b11111111111111;
	assign font[14][252] = 14'b11111111111111;
	assign font[15][252] = 14'b11111111111111;
	assign font[16][252] = 14'b11111111111111;
	assign font[17][252] = 14'b11111111111111;
	assign font[18][252] = 14'b11111111111111;
	assign font[19][252] = 14'b11111111111111;
	assign font[20][252] = 14'b11111111111111;
	assign font[21][252] = 14'b11111111111111;
	assign font[22][252] = 14'b11111111111111;
	assign font[23][252] = 14'b11111111111111;
	assign font[24][252] = 14'b11111111111111;
	assign font[25][252] = 14'b11111111111111;
	assign font[26][252] = 14'b11111111111111;
	assign font[27][252] = 14'b11111111111111;
	assign font[28][252] = 14'b11111111111111;
	assign font[29][252] = 14'b11111111111111;
	assign font[30][252] = 14'b11111111111111;
	assign font[31][252] = 14'b11111111111111;

	assign font[0][253] = 14'b11111111111111;
	assign font[1][253] = 14'b11111111111111;
	assign font[2][253] = 14'b11111111111111;
	assign font[3][253] = 14'b11111111111111;
	assign font[4][253] = 14'b11111111111111;
	assign font[5][253] = 14'b11111111111111;
	assign font[6][253] = 14'b11111111111111;
	assign font[7][253] = 14'b11111111111111;
	assign font[8][253] = 14'b11111111111111;
	assign font[9][253] = 14'b11111111111111;
	assign font[10][253] = 14'b11111111111111;
	assign font[11][253] = 14'b11111111111111;
	assign font[12][253] = 14'b11111111111111;
	assign font[13][253] = 14'b11111111111111;
	assign font[14][253] = 14'b11111111111111;
	assign font[15][253] = 14'b11111111111111;
	assign font[16][253] = 14'b11111111111111;
	assign font[17][253] = 14'b11111111111111;
	assign font[18][253] = 14'b11111111111111;
	assign font[19][253] = 14'b11111111111111;
	assign font[20][253] = 14'b11111111111111;
	assign font[21][253] = 14'b11111111111111;
	assign font[22][253] = 14'b11111111111111;
	assign font[23][253] = 14'b11111111111111;
	assign font[24][253] = 14'b11111111111111;
	assign font[25][253] = 14'b11111111111111;
	assign font[26][253] = 14'b11111111111111;
	assign font[27][253] = 14'b11111111111111;
	assign font[28][253] = 14'b11111111111111;
	assign font[29][253] = 14'b11111111111111;
	assign font[30][253] = 14'b11111111111111;
	assign font[31][253] = 14'b11111111111111;

	assign font[0][254] = 14'b11111111111111;
	assign font[1][254] = 14'b11111111111111;
	assign font[2][254] = 14'b11111111111111;
	assign font[3][254] = 14'b11111111111111;
	assign font[4][254] = 14'b11111111111111;
	assign font[5][254] = 14'b11111111111111;
	assign font[6][254] = 14'b11111111111111;
	assign font[7][254] = 14'b11111111111111;
	assign font[8][254] = 14'b11111111111111;
	assign font[9][254] = 14'b11111111111111;
	assign font[10][254] = 14'b11111111111111;
	assign font[11][254] = 14'b11111111111111;
	assign font[12][254] = 14'b11111111111111;
	assign font[13][254] = 14'b11111111111111;
	assign font[14][254] = 14'b11111111111111;
	assign font[15][254] = 14'b11111111111111;
	assign font[16][254] = 14'b11111111111111;
	assign font[17][254] = 14'b11111111111111;
	assign font[18][254] = 14'b11111111111111;
	assign font[19][254] = 14'b11111111111111;
	assign font[20][254] = 14'b11111111111111;
	assign font[21][254] = 14'b11111111111111;
	assign font[22][254] = 14'b11111111111111;
	assign font[23][254] = 14'b11111111111111;
	assign font[24][254] = 14'b11111111111111;
	assign font[25][254] = 14'b11111111111111;
	assign font[26][254] = 14'b11111111111111;
	assign font[27][254] = 14'b11111111111111;
	assign font[28][254] = 14'b11111111111111;
	assign font[29][254] = 14'b11111111111111;
	assign font[30][254] = 14'b11111111111111;
	assign font[31][254] = 14'b11111111111111;

	assign font[0][255] = 14'b11111111111111;
	assign font[1][255] = 14'b11111111111111;
	assign font[2][255] = 14'b11111111111111;
	assign font[3][255] = 14'b11111111111111;
	assign font[4][255] = 14'b11111111111111;
	assign font[5][255] = 14'b11111111111111;
	assign font[6][255] = 14'b11111111111111;
	assign font[7][255] = 14'b11111111111111;
	assign font[8][255] = 14'b11111111111111;
	assign font[9][255] = 14'b11111111111111;
	assign font[10][255] = 14'b11111111111111;
	assign font[11][255] = 14'b11111111111111;
	assign font[12][255] = 14'b11111111111111;
	assign font[13][255] = 14'b11111111111111;
	assign font[14][255] = 14'b11111111111111;
	assign font[15][255] = 14'b11111111111111;
	assign font[16][255] = 14'b11111111111111;
	assign font[17][255] = 14'b11111111111111;
	assign font[18][255] = 14'b11111111111111;
	assign font[19][255] = 14'b11111111111111;
	assign font[20][255] = 14'b11111111111111;
	assign font[21][255] = 14'b11111111111111;
	assign font[22][255] = 14'b11111111111111;
	assign font[23][255] = 14'b11111111111111;
	assign font[24][255] = 14'b11111111111111;
	assign font[25][255] = 14'b11111111111111;
	assign font[26][255] = 14'b11111111111111;
	assign font[27][255] = 14'b11111111111111;
	assign font[28][255] = 14'b11111111111111;
	assign font[29][255] = 14'b11111111111111;
	assign font[30][255] = 14'b11111111111111;
	assign font[31][255] = 14'b11111111111111;



  assign sym_pixel = font[sym_y][sym_code][sym_x];
endmodule
